module Gowin_DPB (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [31:0] douta;
output [31:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [14:0] ada;
input [31:0] dina;
input [14:0] adb;
input [31:0] dinb;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire [8:0] dpx9b_inst_0_douta_w;
wire [8:0] dpx9b_inst_0_douta;
wire [8:0] dpx9b_inst_0_doutb_w;
wire [8:0] dpx9b_inst_0_doutb;
wire [8:0] dpx9b_inst_1_douta_w;
wire [8:0] dpx9b_inst_1_douta;
wire [8:0] dpx9b_inst_1_doutb_w;
wire [8:0] dpx9b_inst_1_doutb;
wire [8:0] dpx9b_inst_2_douta_w;
wire [8:0] dpx9b_inst_2_douta;
wire [8:0] dpx9b_inst_2_doutb_w;
wire [8:0] dpx9b_inst_2_doutb;
wire [8:0] dpx9b_inst_3_douta_w;
wire [8:0] dpx9b_inst_3_douta;
wire [8:0] dpx9b_inst_3_doutb_w;
wire [8:0] dpx9b_inst_3_doutb;
wire [8:0] dpx9b_inst_4_douta_w;
wire [8:0] dpx9b_inst_4_douta;
wire [8:0] dpx9b_inst_4_doutb_w;
wire [8:0] dpx9b_inst_4_doutb;
wire [8:0] dpx9b_inst_5_douta_w;
wire [8:0] dpx9b_inst_5_douta;
wire [8:0] dpx9b_inst_5_doutb_w;
wire [8:0] dpx9b_inst_5_doutb;
wire [8:0] dpx9b_inst_6_douta_w;
wire [8:0] dpx9b_inst_6_douta;
wire [8:0] dpx9b_inst_6_doutb_w;
wire [8:0] dpx9b_inst_6_doutb;
wire [8:0] dpx9b_inst_7_douta_w;
wire [8:0] dpx9b_inst_7_douta;
wire [8:0] dpx9b_inst_7_doutb_w;
wire [8:0] dpx9b_inst_7_doutb;
wire [8:0] dpx9b_inst_8_douta_w;
wire [8:0] dpx9b_inst_8_douta;
wire [8:0] dpx9b_inst_8_doutb_w;
wire [8:0] dpx9b_inst_8_doutb;
wire [8:0] dpx9b_inst_9_douta_w;
wire [8:0] dpx9b_inst_9_douta;
wire [8:0] dpx9b_inst_9_doutb_w;
wire [8:0] dpx9b_inst_9_doutb;
wire [8:0] dpx9b_inst_10_douta_w;
wire [8:0] dpx9b_inst_10_douta;
wire [8:0] dpx9b_inst_10_doutb_w;
wire [8:0] dpx9b_inst_10_doutb;
wire [8:0] dpx9b_inst_11_douta_w;
wire [8:0] dpx9b_inst_11_douta;
wire [8:0] dpx9b_inst_11_doutb_w;
wire [8:0] dpx9b_inst_11_doutb;
wire [8:0] dpx9b_inst_12_douta_w;
wire [8:0] dpx9b_inst_12_douta;
wire [8:0] dpx9b_inst_12_doutb_w;
wire [8:0] dpx9b_inst_12_doutb;
wire [8:0] dpx9b_inst_13_douta_w;
wire [8:0] dpx9b_inst_13_douta;
wire [8:0] dpx9b_inst_13_doutb_w;
wire [8:0] dpx9b_inst_13_doutb;
wire [8:0] dpx9b_inst_14_douta_w;
wire [17:9] dpx9b_inst_14_douta;
wire [8:0] dpx9b_inst_14_doutb_w;
wire [17:9] dpx9b_inst_14_doutb;
wire [8:0] dpx9b_inst_15_douta_w;
wire [17:9] dpx9b_inst_15_douta;
wire [8:0] dpx9b_inst_15_doutb_w;
wire [17:9] dpx9b_inst_15_doutb;
wire [8:0] dpx9b_inst_16_douta_w;
wire [17:9] dpx9b_inst_16_douta;
wire [8:0] dpx9b_inst_16_doutb_w;
wire [17:9] dpx9b_inst_16_doutb;
wire [8:0] dpx9b_inst_17_douta_w;
wire [17:9] dpx9b_inst_17_douta;
wire [8:0] dpx9b_inst_17_doutb_w;
wire [17:9] dpx9b_inst_17_doutb;
wire [8:0] dpx9b_inst_18_douta_w;
wire [17:9] dpx9b_inst_18_douta;
wire [8:0] dpx9b_inst_18_doutb_w;
wire [17:9] dpx9b_inst_18_doutb;
wire [8:0] dpx9b_inst_19_douta_w;
wire [17:9] dpx9b_inst_19_douta;
wire [8:0] dpx9b_inst_19_doutb_w;
wire [17:9] dpx9b_inst_19_doutb;
wire [8:0] dpx9b_inst_20_douta_w;
wire [17:9] dpx9b_inst_20_douta;
wire [8:0] dpx9b_inst_20_doutb_w;
wire [17:9] dpx9b_inst_20_doutb;
wire [8:0] dpx9b_inst_21_douta_w;
wire [17:9] dpx9b_inst_21_douta;
wire [8:0] dpx9b_inst_21_doutb_w;
wire [17:9] dpx9b_inst_21_doutb;
wire [8:0] dpx9b_inst_22_douta_w;
wire [17:9] dpx9b_inst_22_douta;
wire [8:0] dpx9b_inst_22_doutb_w;
wire [17:9] dpx9b_inst_22_doutb;
wire [8:0] dpx9b_inst_23_douta_w;
wire [17:9] dpx9b_inst_23_douta;
wire [8:0] dpx9b_inst_23_doutb_w;
wire [17:9] dpx9b_inst_23_doutb;
wire [8:0] dpx9b_inst_24_douta_w;
wire [17:9] dpx9b_inst_24_douta;
wire [8:0] dpx9b_inst_24_doutb_w;
wire [17:9] dpx9b_inst_24_doutb;
wire [8:0] dpx9b_inst_25_douta_w;
wire [17:9] dpx9b_inst_25_douta;
wire [8:0] dpx9b_inst_25_doutb_w;
wire [17:9] dpx9b_inst_25_doutb;
wire [8:0] dpx9b_inst_26_douta_w;
wire [17:9] dpx9b_inst_26_douta;
wire [8:0] dpx9b_inst_26_doutb_w;
wire [17:9] dpx9b_inst_26_doutb;
wire [8:0] dpx9b_inst_27_douta_w;
wire [17:9] dpx9b_inst_27_douta;
wire [8:0] dpx9b_inst_27_doutb_w;
wire [17:9] dpx9b_inst_27_doutb;
wire [8:0] dpx9b_inst_28_douta_w;
wire [26:18] dpx9b_inst_28_douta;
wire [8:0] dpx9b_inst_28_doutb_w;
wire [26:18] dpx9b_inst_28_doutb;
wire [8:0] dpx9b_inst_29_douta_w;
wire [26:18] dpx9b_inst_29_douta;
wire [8:0] dpx9b_inst_29_doutb_w;
wire [26:18] dpx9b_inst_29_doutb;
wire [8:0] dpx9b_inst_30_douta_w;
wire [26:18] dpx9b_inst_30_douta;
wire [8:0] dpx9b_inst_30_doutb_w;
wire [26:18] dpx9b_inst_30_doutb;
wire [8:0] dpx9b_inst_31_douta_w;
wire [26:18] dpx9b_inst_31_douta;
wire [8:0] dpx9b_inst_31_doutb_w;
wire [26:18] dpx9b_inst_31_doutb;
wire [8:0] dpx9b_inst_32_douta_w;
wire [26:18] dpx9b_inst_32_douta;
wire [8:0] dpx9b_inst_32_doutb_w;
wire [26:18] dpx9b_inst_32_doutb;
wire [8:0] dpx9b_inst_33_douta_w;
wire [26:18] dpx9b_inst_33_douta;
wire [8:0] dpx9b_inst_33_doutb_w;
wire [26:18] dpx9b_inst_33_doutb;
wire [8:0] dpx9b_inst_34_douta_w;
wire [26:18] dpx9b_inst_34_douta;
wire [8:0] dpx9b_inst_34_doutb_w;
wire [26:18] dpx9b_inst_34_doutb;
wire [8:0] dpx9b_inst_35_douta_w;
wire [26:18] dpx9b_inst_35_douta;
wire [8:0] dpx9b_inst_35_doutb_w;
wire [26:18] dpx9b_inst_35_doutb;
wire [8:0] dpx9b_inst_36_douta_w;
wire [26:18] dpx9b_inst_36_douta;
wire [8:0] dpx9b_inst_36_doutb_w;
wire [26:18] dpx9b_inst_36_doutb;
wire [8:0] dpx9b_inst_37_douta_w;
wire [26:18] dpx9b_inst_37_douta;
wire [8:0] dpx9b_inst_37_doutb_w;
wire [26:18] dpx9b_inst_37_doutb;
wire [8:0] dpx9b_inst_38_douta_w;
wire [26:18] dpx9b_inst_38_douta;
wire [8:0] dpx9b_inst_38_doutb_w;
wire [26:18] dpx9b_inst_38_doutb;
wire [8:0] dpx9b_inst_39_douta_w;
wire [26:18] dpx9b_inst_39_douta;
wire [8:0] dpx9b_inst_39_doutb_w;
wire [26:18] dpx9b_inst_39_doutb;
wire [8:0] dpx9b_inst_40_douta_w;
wire [26:18] dpx9b_inst_40_douta;
wire [8:0] dpx9b_inst_40_doutb_w;
wire [26:18] dpx9b_inst_40_doutb;
wire [8:0] dpx9b_inst_41_douta_w;
wire [26:18] dpx9b_inst_41_douta;
wire [8:0] dpx9b_inst_41_doutb_w;
wire [26:18] dpx9b_inst_41_doutb;
wire [14:0] dpb_inst_42_douta_w;
wire [27:27] dpb_inst_42_douta;
wire [14:0] dpb_inst_42_doutb_w;
wire [27:27] dpb_inst_42_doutb;
wire [14:0] dpb_inst_43_douta_w;
wire [28:28] dpb_inst_43_douta;
wire [14:0] dpb_inst_43_doutb_w;
wire [28:28] dpb_inst_43_doutb;
wire [14:0] dpb_inst_44_douta_w;
wire [29:29] dpb_inst_44_douta;
wire [14:0] dpb_inst_44_doutb_w;
wire [29:29] dpb_inst_44_doutb;
wire [14:0] dpb_inst_45_douta_w;
wire [30:30] dpb_inst_45_douta;
wire [14:0] dpb_inst_45_doutb_w;
wire [30:30] dpb_inst_45_doutb;
wire [13:0] dpb_inst_46_douta_w;
wire [28:27] dpb_inst_46_douta;
wire [13:0] dpb_inst_46_doutb_w;
wire [28:27] dpb_inst_46_doutb;
wire [13:0] dpb_inst_47_douta_w;
wire [30:29] dpb_inst_47_douta;
wire [13:0] dpb_inst_47_doutb_w;
wire [30:29] dpb_inst_47_doutb;
wire [11:0] dpb_inst_48_douta_w;
wire [30:27] dpb_inst_48_douta;
wire [11:0] dpb_inst_48_doutb_w;
wire [30:27] dpb_inst_48_doutb;
wire [14:0] dpb_inst_49_douta_w;
wire [31:31] dpb_inst_49_douta;
wire [14:0] dpb_inst_49_doutb_w;
wire [31:31] dpb_inst_49_doutb;
wire [14:0] dpb_inst_50_douta_w;
wire [31:31] dpb_inst_50_douta;
wire [14:0] dpb_inst_50_doutb_w;
wire [31:31] dpb_inst_50_doutb;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire dff_q_6;
wire dff_q_7;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_11;
wire mux_o_12;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_25;
wire mux_o_26;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_39;
wire mux_o_40;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_53;
wire mux_o_54;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_67;
wire mux_o_68;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_81;
wire mux_o_82;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_95;
wire mux_o_96;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_104;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_109;
wire mux_o_110;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_123;
wire mux_o_124;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_137;
wire mux_o_138;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_151;
wire mux_o_152;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_165;
wire mux_o_166;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_179;
wire mux_o_180;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_193;
wire mux_o_194;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_207;
wire mux_o_208;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_221;
wire mux_o_222;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_235;
wire mux_o_236;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_249;
wire mux_o_250;
wire mux_o_252;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_263;
wire mux_o_264;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_277;
wire mux_o_278;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_291;
wire mux_o_292;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_305;
wire mux_o_306;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_314;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_319;
wire mux_o_320;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_333;
wire mux_o_334;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_347;
wire mux_o_348;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_361;
wire mux_o_362;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_375;
wire mux_o_376;
wire mux_o_385;
wire mux_o_394;
wire mux_o_403;
wire mux_o_412;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_432;
wire mux_o_433;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_440;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_446;
wire mux_o_447;
wire mux_o_449;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_460;
wire mux_o_461;
wire mux_o_463;
wire mux_o_464;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_474;
wire mux_o_475;
wire mux_o_477;
wire mux_o_478;
wire mux_o_479;
wire mux_o_480;
wire mux_o_481;
wire mux_o_482;
wire mux_o_483;
wire mux_o_484;
wire mux_o_485;
wire mux_o_486;
wire mux_o_488;
wire mux_o_489;
wire mux_o_491;
wire mux_o_492;
wire mux_o_493;
wire mux_o_494;
wire mux_o_495;
wire mux_o_496;
wire mux_o_497;
wire mux_o_498;
wire mux_o_499;
wire mux_o_500;
wire mux_o_502;
wire mux_o_503;
wire mux_o_505;
wire mux_o_506;
wire mux_o_507;
wire mux_o_508;
wire mux_o_509;
wire mux_o_510;
wire mux_o_511;
wire mux_o_512;
wire mux_o_513;
wire mux_o_514;
wire mux_o_516;
wire mux_o_517;
wire mux_o_519;
wire mux_o_520;
wire mux_o_521;
wire mux_o_522;
wire mux_o_523;
wire mux_o_524;
wire mux_o_525;
wire mux_o_526;
wire mux_o_527;
wire mux_o_528;
wire mux_o_530;
wire mux_o_531;
wire mux_o_533;
wire mux_o_534;
wire mux_o_535;
wire mux_o_536;
wire mux_o_537;
wire mux_o_538;
wire mux_o_539;
wire mux_o_540;
wire mux_o_541;
wire mux_o_542;
wire mux_o_544;
wire mux_o_545;
wire mux_o_547;
wire mux_o_548;
wire mux_o_549;
wire mux_o_550;
wire mux_o_551;
wire mux_o_552;
wire mux_o_553;
wire mux_o_554;
wire mux_o_555;
wire mux_o_556;
wire mux_o_558;
wire mux_o_559;
wire mux_o_561;
wire mux_o_562;
wire mux_o_563;
wire mux_o_564;
wire mux_o_565;
wire mux_o_566;
wire mux_o_567;
wire mux_o_568;
wire mux_o_569;
wire mux_o_570;
wire mux_o_572;
wire mux_o_573;
wire mux_o_575;
wire mux_o_576;
wire mux_o_577;
wire mux_o_578;
wire mux_o_579;
wire mux_o_580;
wire mux_o_581;
wire mux_o_582;
wire mux_o_583;
wire mux_o_584;
wire mux_o_586;
wire mux_o_587;
wire mux_o_589;
wire mux_o_590;
wire mux_o_591;
wire mux_o_592;
wire mux_o_593;
wire mux_o_594;
wire mux_o_595;
wire mux_o_596;
wire mux_o_597;
wire mux_o_598;
wire mux_o_600;
wire mux_o_601;
wire mux_o_603;
wire mux_o_604;
wire mux_o_605;
wire mux_o_606;
wire mux_o_607;
wire mux_o_608;
wire mux_o_609;
wire mux_o_610;
wire mux_o_611;
wire mux_o_612;
wire mux_o_614;
wire mux_o_615;
wire mux_o_617;
wire mux_o_618;
wire mux_o_619;
wire mux_o_620;
wire mux_o_621;
wire mux_o_622;
wire mux_o_623;
wire mux_o_624;
wire mux_o_625;
wire mux_o_626;
wire mux_o_628;
wire mux_o_629;
wire mux_o_631;
wire mux_o_632;
wire mux_o_633;
wire mux_o_634;
wire mux_o_635;
wire mux_o_636;
wire mux_o_637;
wire mux_o_638;
wire mux_o_639;
wire mux_o_640;
wire mux_o_642;
wire mux_o_643;
wire mux_o_645;
wire mux_o_646;
wire mux_o_647;
wire mux_o_648;
wire mux_o_649;
wire mux_o_650;
wire mux_o_651;
wire mux_o_652;
wire mux_o_653;
wire mux_o_654;
wire mux_o_656;
wire mux_o_657;
wire mux_o_659;
wire mux_o_660;
wire mux_o_661;
wire mux_o_662;
wire mux_o_663;
wire mux_o_664;
wire mux_o_665;
wire mux_o_666;
wire mux_o_667;
wire mux_o_668;
wire mux_o_670;
wire mux_o_671;
wire mux_o_673;
wire mux_o_674;
wire mux_o_675;
wire mux_o_676;
wire mux_o_677;
wire mux_o_678;
wire mux_o_679;
wire mux_o_680;
wire mux_o_681;
wire mux_o_682;
wire mux_o_684;
wire mux_o_685;
wire mux_o_687;
wire mux_o_688;
wire mux_o_689;
wire mux_o_690;
wire mux_o_691;
wire mux_o_692;
wire mux_o_693;
wire mux_o_694;
wire mux_o_695;
wire mux_o_696;
wire mux_o_698;
wire mux_o_699;
wire mux_o_701;
wire mux_o_702;
wire mux_o_703;
wire mux_o_704;
wire mux_o_705;
wire mux_o_706;
wire mux_o_707;
wire mux_o_708;
wire mux_o_709;
wire mux_o_710;
wire mux_o_712;
wire mux_o_713;
wire mux_o_715;
wire mux_o_716;
wire mux_o_717;
wire mux_o_718;
wire mux_o_719;
wire mux_o_720;
wire mux_o_721;
wire mux_o_722;
wire mux_o_723;
wire mux_o_724;
wire mux_o_726;
wire mux_o_727;
wire mux_o_729;
wire mux_o_730;
wire mux_o_731;
wire mux_o_732;
wire mux_o_733;
wire mux_o_734;
wire mux_o_735;
wire mux_o_736;
wire mux_o_737;
wire mux_o_738;
wire mux_o_740;
wire mux_o_741;
wire mux_o_743;
wire mux_o_744;
wire mux_o_745;
wire mux_o_746;
wire mux_o_747;
wire mux_o_748;
wire mux_o_749;
wire mux_o_750;
wire mux_o_751;
wire mux_o_752;
wire mux_o_754;
wire mux_o_755;
wire mux_o_757;
wire mux_o_758;
wire mux_o_759;
wire mux_o_760;
wire mux_o_761;
wire mux_o_762;
wire mux_o_763;
wire mux_o_764;
wire mux_o_765;
wire mux_o_766;
wire mux_o_768;
wire mux_o_769;
wire mux_o_771;
wire mux_o_772;
wire mux_o_773;
wire mux_o_774;
wire mux_o_775;
wire mux_o_776;
wire mux_o_777;
wire mux_o_778;
wire mux_o_779;
wire mux_o_780;
wire mux_o_782;
wire mux_o_783;
wire mux_o_785;
wire mux_o_786;
wire mux_o_787;
wire mux_o_788;
wire mux_o_789;
wire mux_o_790;
wire mux_o_791;
wire mux_o_792;
wire mux_o_793;
wire mux_o_794;
wire mux_o_796;
wire mux_o_797;
wire mux_o_806;
wire mux_o_815;
wire mux_o_824;
wire mux_o_833;
wire cea_w;
wire ceb_w;
wire gw_gnd;

assign cea_w = ~wrea & cea;
assign ceb_w = ~wreb & ceb;
assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_0.INIT = 16'h0001;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_1.INIT = 16'h0002;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_2.INIT = 16'h0004;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_3.INIT = 16'h0008;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_4.INIT = 16'h0010;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_5.INIT = 16'h0020;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_6.INIT = 16'h0040;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_7.INIT = 16'h0080;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_8.INIT = 16'h0100;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_9.INIT = 16'h0200;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_10.INIT = 16'h0400;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_11.INIT = 16'h0800;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_12.INIT = 16'h1000;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_13.INIT = 16'h2000;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_14.INIT = 16'h0001;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_15.INIT = 16'h0002;
LUT4 lut_inst_16 (
  .F(lut_f_16),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_16.INIT = 16'h0004;
LUT4 lut_inst_17 (
  .F(lut_f_17),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_17.INIT = 16'h0008;
LUT4 lut_inst_18 (
  .F(lut_f_18),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_18.INIT = 16'h0010;
LUT4 lut_inst_19 (
  .F(lut_f_19),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_19.INIT = 16'h0020;
LUT4 lut_inst_20 (
  .F(lut_f_20),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_20.INIT = 16'h0040;
LUT4 lut_inst_21 (
  .F(lut_f_21),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_21.INIT = 16'h0080;
LUT4 lut_inst_22 (
  .F(lut_f_22),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_22.INIT = 16'h0100;
LUT4 lut_inst_23 (
  .F(lut_f_23),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_23.INIT = 16'h0200;
LUT4 lut_inst_24 (
  .F(lut_f_24),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_24.INIT = 16'h0400;
LUT4 lut_inst_25 (
  .F(lut_f_25),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_25.INIT = 16'h0800;
LUT4 lut_inst_26 (
  .F(lut_f_26),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_26.INIT = 16'h1000;
LUT4 lut_inst_27 (
  .F(lut_f_27),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_27.INIT = 16'h2000;
DPX9B dpx9b_inst_0 (
    .DOA({dpx9b_inst_0_douta_w[8:0],dpx9b_inst_0_douta[8:0]}),
    .DOB({dpx9b_inst_0_doutb_w[8:0],dpx9b_inst_0_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_14}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_0.READ_MODE0 = 1'b0;
defparam dpx9b_inst_0.READ_MODE1 = 1'b0;
defparam dpx9b_inst_0.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_0.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_0.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_0.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_0.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_0.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_0.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_1 (
    .DOA({dpx9b_inst_1_douta_w[8:0],dpx9b_inst_1_douta[8:0]}),
    .DOB({dpx9b_inst_1_doutb_w[8:0],dpx9b_inst_1_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_15}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_1.READ_MODE0 = 1'b0;
defparam dpx9b_inst_1.READ_MODE1 = 1'b0;
defparam dpx9b_inst_1.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_1.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_1.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_1.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_1.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_1.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_1.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_2 (
    .DOA({dpx9b_inst_2_douta_w[8:0],dpx9b_inst_2_douta[8:0]}),
    .DOB({dpx9b_inst_2_doutb_w[8:0],dpx9b_inst_2_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_16}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_2.READ_MODE0 = 1'b0;
defparam dpx9b_inst_2.READ_MODE1 = 1'b0;
defparam dpx9b_inst_2.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_2.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_2.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_2.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_2.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_2.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_2.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_3 (
    .DOA({dpx9b_inst_3_douta_w[8:0],dpx9b_inst_3_douta[8:0]}),
    .DOB({dpx9b_inst_3_doutb_w[8:0],dpx9b_inst_3_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_17}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_3.READ_MODE0 = 1'b0;
defparam dpx9b_inst_3.READ_MODE1 = 1'b0;
defparam dpx9b_inst_3.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_3.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_3.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_3.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_3.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_3.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_3.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_4 (
    .DOA({dpx9b_inst_4_douta_w[8:0],dpx9b_inst_4_douta[8:0]}),
    .DOB({dpx9b_inst_4_doutb_w[8:0],dpx9b_inst_4_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_18}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_4.READ_MODE0 = 1'b0;
defparam dpx9b_inst_4.READ_MODE1 = 1'b0;
defparam dpx9b_inst_4.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_4.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_4.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_4.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_4.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_4.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_4.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_5 (
    .DOA({dpx9b_inst_5_douta_w[8:0],dpx9b_inst_5_douta[8:0]}),
    .DOB({dpx9b_inst_5_doutb_w[8:0],dpx9b_inst_5_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_19}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_5.READ_MODE0 = 1'b0;
defparam dpx9b_inst_5.READ_MODE1 = 1'b0;
defparam dpx9b_inst_5.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_5.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_5.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_5.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_5.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_5.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_5.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_6 (
    .DOA({dpx9b_inst_6_douta_w[8:0],dpx9b_inst_6_douta[8:0]}),
    .DOB({dpx9b_inst_6_doutb_w[8:0],dpx9b_inst_6_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_20}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_6.READ_MODE0 = 1'b0;
defparam dpx9b_inst_6.READ_MODE1 = 1'b0;
defparam dpx9b_inst_6.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_6.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_6.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_6.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_6.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_6.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_6.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_7 (
    .DOA({dpx9b_inst_7_douta_w[8:0],dpx9b_inst_7_douta[8:0]}),
    .DOB({dpx9b_inst_7_doutb_w[8:0],dpx9b_inst_7_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_21}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_7.READ_MODE0 = 1'b0;
defparam dpx9b_inst_7.READ_MODE1 = 1'b0;
defparam dpx9b_inst_7.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_7.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_7.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_7.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_7.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_7.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_7.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_8 (
    .DOA({dpx9b_inst_8_douta_w[8:0],dpx9b_inst_8_douta[8:0]}),
    .DOB({dpx9b_inst_8_doutb_w[8:0],dpx9b_inst_8_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_22}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_8.READ_MODE0 = 1'b0;
defparam dpx9b_inst_8.READ_MODE1 = 1'b0;
defparam dpx9b_inst_8.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_8.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_8.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_8.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_8.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_8.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_8.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_9 (
    .DOA({dpx9b_inst_9_douta_w[8:0],dpx9b_inst_9_douta[8:0]}),
    .DOB({dpx9b_inst_9_doutb_w[8:0],dpx9b_inst_9_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_23}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_9.READ_MODE0 = 1'b0;
defparam dpx9b_inst_9.READ_MODE1 = 1'b0;
defparam dpx9b_inst_9.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_9.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_9.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_9.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_9.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_9.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_9.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_10 (
    .DOA({dpx9b_inst_10_douta_w[8:0],dpx9b_inst_10_douta[8:0]}),
    .DOB({dpx9b_inst_10_doutb_w[8:0],dpx9b_inst_10_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_24}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_10.READ_MODE0 = 1'b0;
defparam dpx9b_inst_10.READ_MODE1 = 1'b0;
defparam dpx9b_inst_10.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_10.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_10.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_10.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_10.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_10.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_10.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_11 (
    .DOA({dpx9b_inst_11_douta_w[8:0],dpx9b_inst_11_douta[8:0]}),
    .DOB({dpx9b_inst_11_doutb_w[8:0],dpx9b_inst_11_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_25}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_11.READ_MODE0 = 1'b0;
defparam dpx9b_inst_11.READ_MODE1 = 1'b0;
defparam dpx9b_inst_11.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_11.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_11.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_11.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_11.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_11.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_11.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_12 (
    .DOA({dpx9b_inst_12_douta_w[8:0],dpx9b_inst_12_douta[8:0]}),
    .DOB({dpx9b_inst_12_doutb_w[8:0],dpx9b_inst_12_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_26}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_12.READ_MODE0 = 1'b0;
defparam dpx9b_inst_12.READ_MODE1 = 1'b0;
defparam dpx9b_inst_12.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_12.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_12.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_12.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_12.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_12.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_12.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_13 (
    .DOA({dpx9b_inst_13_douta_w[8:0],dpx9b_inst_13_douta[8:0]}),
    .DOB({dpx9b_inst_13_doutb_w[8:0],dpx9b_inst_13_doutb[8:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_27}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[8:0]})
);

defparam dpx9b_inst_13.READ_MODE0 = 1'b0;
defparam dpx9b_inst_13.READ_MODE1 = 1'b0;
defparam dpx9b_inst_13.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_13.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_13.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_13.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_13.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_13.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_13.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_14 (
    .DOA({dpx9b_inst_14_douta_w[8:0],dpx9b_inst_14_douta[17:9]}),
    .DOB({dpx9b_inst_14_doutb_w[8:0],dpx9b_inst_14_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_14}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_14.READ_MODE0 = 1'b0;
defparam dpx9b_inst_14.READ_MODE1 = 1'b0;
defparam dpx9b_inst_14.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_14.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_14.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_14.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_14.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_14.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_14.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_15 (
    .DOA({dpx9b_inst_15_douta_w[8:0],dpx9b_inst_15_douta[17:9]}),
    .DOB({dpx9b_inst_15_doutb_w[8:0],dpx9b_inst_15_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_15}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_15.READ_MODE0 = 1'b0;
defparam dpx9b_inst_15.READ_MODE1 = 1'b0;
defparam dpx9b_inst_15.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_15.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_15.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_15.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_15.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_15.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_15.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_16 (
    .DOA({dpx9b_inst_16_douta_w[8:0],dpx9b_inst_16_douta[17:9]}),
    .DOB({dpx9b_inst_16_doutb_w[8:0],dpx9b_inst_16_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_16}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_16.READ_MODE0 = 1'b0;
defparam dpx9b_inst_16.READ_MODE1 = 1'b0;
defparam dpx9b_inst_16.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_16.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_16.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_16.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_16.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_16.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_16.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_17 (
    .DOA({dpx9b_inst_17_douta_w[8:0],dpx9b_inst_17_douta[17:9]}),
    .DOB({dpx9b_inst_17_doutb_w[8:0],dpx9b_inst_17_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_17}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_17.READ_MODE0 = 1'b0;
defparam dpx9b_inst_17.READ_MODE1 = 1'b0;
defparam dpx9b_inst_17.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_17.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_17.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_17.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_17.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_17.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_17.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_18 (
    .DOA({dpx9b_inst_18_douta_w[8:0],dpx9b_inst_18_douta[17:9]}),
    .DOB({dpx9b_inst_18_doutb_w[8:0],dpx9b_inst_18_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_18}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_18.READ_MODE0 = 1'b0;
defparam dpx9b_inst_18.READ_MODE1 = 1'b0;
defparam dpx9b_inst_18.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_18.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_18.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_18.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_18.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_18.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_18.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_19 (
    .DOA({dpx9b_inst_19_douta_w[8:0],dpx9b_inst_19_douta[17:9]}),
    .DOB({dpx9b_inst_19_doutb_w[8:0],dpx9b_inst_19_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_19}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_19.READ_MODE0 = 1'b0;
defparam dpx9b_inst_19.READ_MODE1 = 1'b0;
defparam dpx9b_inst_19.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_19.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_19.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_19.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_19.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_19.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_19.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_20 (
    .DOA({dpx9b_inst_20_douta_w[8:0],dpx9b_inst_20_douta[17:9]}),
    .DOB({dpx9b_inst_20_doutb_w[8:0],dpx9b_inst_20_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_20}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_20.READ_MODE0 = 1'b0;
defparam dpx9b_inst_20.READ_MODE1 = 1'b0;
defparam dpx9b_inst_20.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_20.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_20.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_20.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_20.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_20.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_20.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_21 (
    .DOA({dpx9b_inst_21_douta_w[8:0],dpx9b_inst_21_douta[17:9]}),
    .DOB({dpx9b_inst_21_doutb_w[8:0],dpx9b_inst_21_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_21}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_21.READ_MODE0 = 1'b0;
defparam dpx9b_inst_21.READ_MODE1 = 1'b0;
defparam dpx9b_inst_21.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_21.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_21.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_21.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_21.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_21.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_21.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_22 (
    .DOA({dpx9b_inst_22_douta_w[8:0],dpx9b_inst_22_douta[17:9]}),
    .DOB({dpx9b_inst_22_doutb_w[8:0],dpx9b_inst_22_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_22}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_22.READ_MODE0 = 1'b0;
defparam dpx9b_inst_22.READ_MODE1 = 1'b0;
defparam dpx9b_inst_22.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_22.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_22.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_22.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_22.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_22.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_22.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_23 (
    .DOA({dpx9b_inst_23_douta_w[8:0],dpx9b_inst_23_douta[17:9]}),
    .DOB({dpx9b_inst_23_doutb_w[8:0],dpx9b_inst_23_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_23}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_23.READ_MODE0 = 1'b0;
defparam dpx9b_inst_23.READ_MODE1 = 1'b0;
defparam dpx9b_inst_23.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_23.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_23.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_23.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_23.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_23.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_23.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_24 (
    .DOA({dpx9b_inst_24_douta_w[8:0],dpx9b_inst_24_douta[17:9]}),
    .DOB({dpx9b_inst_24_doutb_w[8:0],dpx9b_inst_24_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_24}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_24.READ_MODE0 = 1'b0;
defparam dpx9b_inst_24.READ_MODE1 = 1'b0;
defparam dpx9b_inst_24.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_24.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_24.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_24.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_24.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_24.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_24.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_25 (
    .DOA({dpx9b_inst_25_douta_w[8:0],dpx9b_inst_25_douta[17:9]}),
    .DOB({dpx9b_inst_25_doutb_w[8:0],dpx9b_inst_25_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_25}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_25.READ_MODE0 = 1'b0;
defparam dpx9b_inst_25.READ_MODE1 = 1'b0;
defparam dpx9b_inst_25.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_25.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_25.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_25.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_25.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_25.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_25.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_26 (
    .DOA({dpx9b_inst_26_douta_w[8:0],dpx9b_inst_26_douta[17:9]}),
    .DOB({dpx9b_inst_26_doutb_w[8:0],dpx9b_inst_26_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_26}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_26.READ_MODE0 = 1'b0;
defparam dpx9b_inst_26.READ_MODE1 = 1'b0;
defparam dpx9b_inst_26.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_26.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_26.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_26.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_26.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_26.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_26.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_27 (
    .DOA({dpx9b_inst_27_douta_w[8:0],dpx9b_inst_27_douta[17:9]}),
    .DOB({dpx9b_inst_27_doutb_w[8:0],dpx9b_inst_27_doutb[17:9]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_27}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[17:9]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[17:9]})
);

defparam dpx9b_inst_27.READ_MODE0 = 1'b0;
defparam dpx9b_inst_27.READ_MODE1 = 1'b0;
defparam dpx9b_inst_27.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_27.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_27.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_27.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_27.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_27.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_27.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_28 (
    .DOA({dpx9b_inst_28_douta_w[8:0],dpx9b_inst_28_douta[26:18]}),
    .DOB({dpx9b_inst_28_doutb_w[8:0],dpx9b_inst_28_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_14}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_28.READ_MODE0 = 1'b0;
defparam dpx9b_inst_28.READ_MODE1 = 1'b0;
defparam dpx9b_inst_28.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_28.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_28.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_28.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_28.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_28.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_28.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_29 (
    .DOA({dpx9b_inst_29_douta_w[8:0],dpx9b_inst_29_douta[26:18]}),
    .DOB({dpx9b_inst_29_doutb_w[8:0],dpx9b_inst_29_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_15}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_29.READ_MODE0 = 1'b0;
defparam dpx9b_inst_29.READ_MODE1 = 1'b0;
defparam dpx9b_inst_29.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_29.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_29.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_29.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_29.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_29.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_29.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_30 (
    .DOA({dpx9b_inst_30_douta_w[8:0],dpx9b_inst_30_douta[26:18]}),
    .DOB({dpx9b_inst_30_doutb_w[8:0],dpx9b_inst_30_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_16}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_30.READ_MODE0 = 1'b0;
defparam dpx9b_inst_30.READ_MODE1 = 1'b0;
defparam dpx9b_inst_30.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_30.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_30.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_30.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_30.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_30.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_30.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_31 (
    .DOA({dpx9b_inst_31_douta_w[8:0],dpx9b_inst_31_douta[26:18]}),
    .DOB({dpx9b_inst_31_doutb_w[8:0],dpx9b_inst_31_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_17}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_31.READ_MODE0 = 1'b0;
defparam dpx9b_inst_31.READ_MODE1 = 1'b0;
defparam dpx9b_inst_31.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_31.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_31.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_31.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_31.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_31.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_31.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_32 (
    .DOA({dpx9b_inst_32_douta_w[8:0],dpx9b_inst_32_douta[26:18]}),
    .DOB({dpx9b_inst_32_doutb_w[8:0],dpx9b_inst_32_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_18}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_32.READ_MODE0 = 1'b0;
defparam dpx9b_inst_32.READ_MODE1 = 1'b0;
defparam dpx9b_inst_32.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_32.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_32.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_32.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_32.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_32.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_32.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_33 (
    .DOA({dpx9b_inst_33_douta_w[8:0],dpx9b_inst_33_douta[26:18]}),
    .DOB({dpx9b_inst_33_doutb_w[8:0],dpx9b_inst_33_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_19}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_33.READ_MODE0 = 1'b0;
defparam dpx9b_inst_33.READ_MODE1 = 1'b0;
defparam dpx9b_inst_33.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_33.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_33.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_33.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_33.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_33.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_33.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_34 (
    .DOA({dpx9b_inst_34_douta_w[8:0],dpx9b_inst_34_douta[26:18]}),
    .DOB({dpx9b_inst_34_doutb_w[8:0],dpx9b_inst_34_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_20}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_34.READ_MODE0 = 1'b0;
defparam dpx9b_inst_34.READ_MODE1 = 1'b0;
defparam dpx9b_inst_34.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_34.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_34.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_34.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_34.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_34.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_34.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_35 (
    .DOA({dpx9b_inst_35_douta_w[8:0],dpx9b_inst_35_douta[26:18]}),
    .DOB({dpx9b_inst_35_doutb_w[8:0],dpx9b_inst_35_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_21}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_35.READ_MODE0 = 1'b0;
defparam dpx9b_inst_35.READ_MODE1 = 1'b0;
defparam dpx9b_inst_35.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_35.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_35.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_35.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_35.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_35.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_35.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_36 (
    .DOA({dpx9b_inst_36_douta_w[8:0],dpx9b_inst_36_douta[26:18]}),
    .DOB({dpx9b_inst_36_doutb_w[8:0],dpx9b_inst_36_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_22}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_36.READ_MODE0 = 1'b0;
defparam dpx9b_inst_36.READ_MODE1 = 1'b0;
defparam dpx9b_inst_36.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_36.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_36.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_36.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_36.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_36.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_36.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_37 (
    .DOA({dpx9b_inst_37_douta_w[8:0],dpx9b_inst_37_douta[26:18]}),
    .DOB({dpx9b_inst_37_doutb_w[8:0],dpx9b_inst_37_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_23}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_37.READ_MODE0 = 1'b0;
defparam dpx9b_inst_37.READ_MODE1 = 1'b0;
defparam dpx9b_inst_37.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_37.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_37.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_37.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_37.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_37.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_37.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_38 (
    .DOA({dpx9b_inst_38_douta_w[8:0],dpx9b_inst_38_douta[26:18]}),
    .DOB({dpx9b_inst_38_doutb_w[8:0],dpx9b_inst_38_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_24}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_38.READ_MODE0 = 1'b0;
defparam dpx9b_inst_38.READ_MODE1 = 1'b0;
defparam dpx9b_inst_38.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_38.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_38.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_38.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_38.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_38.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_38.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_39 (
    .DOA({dpx9b_inst_39_douta_w[8:0],dpx9b_inst_39_douta[26:18]}),
    .DOB({dpx9b_inst_39_doutb_w[8:0],dpx9b_inst_39_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_25}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_39.READ_MODE0 = 1'b0;
defparam dpx9b_inst_39.READ_MODE1 = 1'b0;
defparam dpx9b_inst_39.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_39.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_39.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_39.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_39.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_39.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_39.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_40 (
    .DOA({dpx9b_inst_40_douta_w[8:0],dpx9b_inst_40_douta[26:18]}),
    .DOB({dpx9b_inst_40_doutb_w[8:0],dpx9b_inst_40_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_26}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_40.READ_MODE0 = 1'b0;
defparam dpx9b_inst_40.READ_MODE1 = 1'b0;
defparam dpx9b_inst_40.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_40.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_40.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_40.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_40.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_40.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_40.RESET_MODE = "SYNC";

DPX9B dpx9b_inst_41 (
    .DOA({dpx9b_inst_41_douta_w[8:0],dpx9b_inst_41_douta[26:18]}),
    .DOB({dpx9b_inst_41_doutb_w[8:0],dpx9b_inst_41_doutb[26:18]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_27}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[26:18]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[26:18]})
);

defparam dpx9b_inst_41.READ_MODE0 = 1'b0;
defparam dpx9b_inst_41.READ_MODE1 = 1'b0;
defparam dpx9b_inst_41.WRITE_MODE0 = 2'b00;
defparam dpx9b_inst_41.WRITE_MODE1 = 2'b00;
defparam dpx9b_inst_41.BIT_WIDTH_0 = 9;
defparam dpx9b_inst_41.BIT_WIDTH_1 = 9;
defparam dpx9b_inst_41.BLK_SEL_0 = 3'b001;
defparam dpx9b_inst_41.BLK_SEL_1 = 3'b001;
defparam dpx9b_inst_41.RESET_MODE = "SYNC";

DPB dpb_inst_42 (
    .DOA({dpb_inst_42_douta_w[14:0],dpb_inst_42_douta[27]}),
    .DOB({dpb_inst_42_doutb_w[14:0],dpb_inst_42_doutb[27]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[27]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[27]})
);

defparam dpb_inst_42.READ_MODE0 = 1'b0;
defparam dpb_inst_42.READ_MODE1 = 1'b0;
defparam dpb_inst_42.WRITE_MODE0 = 2'b00;
defparam dpb_inst_42.WRITE_MODE1 = 2'b00;
defparam dpb_inst_42.BIT_WIDTH_0 = 1;
defparam dpb_inst_42.BIT_WIDTH_1 = 1;
defparam dpb_inst_42.BLK_SEL_0 = 3'b000;
defparam dpb_inst_42.BLK_SEL_1 = 3'b000;
defparam dpb_inst_42.RESET_MODE = "SYNC";

DPB dpb_inst_43 (
    .DOA({dpb_inst_43_douta_w[14:0],dpb_inst_43_douta[28]}),
    .DOB({dpb_inst_43_doutb_w[14:0],dpb_inst_43_doutb[28]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[28]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[28]})
);

defparam dpb_inst_43.READ_MODE0 = 1'b0;
defparam dpb_inst_43.READ_MODE1 = 1'b0;
defparam dpb_inst_43.WRITE_MODE0 = 2'b00;
defparam dpb_inst_43.WRITE_MODE1 = 2'b00;
defparam dpb_inst_43.BIT_WIDTH_0 = 1;
defparam dpb_inst_43.BIT_WIDTH_1 = 1;
defparam dpb_inst_43.BLK_SEL_0 = 3'b000;
defparam dpb_inst_43.BLK_SEL_1 = 3'b000;
defparam dpb_inst_43.RESET_MODE = "SYNC";

DPB dpb_inst_44 (
    .DOA({dpb_inst_44_douta_w[14:0],dpb_inst_44_douta[29]}),
    .DOB({dpb_inst_44_doutb_w[14:0],dpb_inst_44_doutb[29]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[29]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[29]})
);

defparam dpb_inst_44.READ_MODE0 = 1'b0;
defparam dpb_inst_44.READ_MODE1 = 1'b0;
defparam dpb_inst_44.WRITE_MODE0 = 2'b00;
defparam dpb_inst_44.WRITE_MODE1 = 2'b00;
defparam dpb_inst_44.BIT_WIDTH_0 = 1;
defparam dpb_inst_44.BIT_WIDTH_1 = 1;
defparam dpb_inst_44.BLK_SEL_0 = 3'b000;
defparam dpb_inst_44.BLK_SEL_1 = 3'b000;
defparam dpb_inst_44.RESET_MODE = "SYNC";

DPB dpb_inst_45 (
    .DOA({dpb_inst_45_douta_w[14:0],dpb_inst_45_douta[30]}),
    .DOB({dpb_inst_45_doutb_w[14:0],dpb_inst_45_doutb[30]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[30]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[30]})
);

defparam dpb_inst_45.READ_MODE0 = 1'b0;
defparam dpb_inst_45.READ_MODE1 = 1'b0;
defparam dpb_inst_45.WRITE_MODE0 = 2'b00;
defparam dpb_inst_45.WRITE_MODE1 = 2'b00;
defparam dpb_inst_45.BIT_WIDTH_0 = 1;
defparam dpb_inst_45.BIT_WIDTH_1 = 1;
defparam dpb_inst_45.BLK_SEL_0 = 3'b000;
defparam dpb_inst_45.BLK_SEL_1 = 3'b000;
defparam dpb_inst_45.RESET_MODE = "SYNC";

DPB dpb_inst_46 (
    .DOA({dpb_inst_46_douta_w[13:0],dpb_inst_46_douta[28:27]}),
    .DOB({dpb_inst_46_doutb_w[13:0],dpb_inst_46_doutb[28:27]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[28:27]}),
    .ADB({adb[12:0],gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[28:27]})
);

defparam dpb_inst_46.READ_MODE0 = 1'b0;
defparam dpb_inst_46.READ_MODE1 = 1'b0;
defparam dpb_inst_46.WRITE_MODE0 = 2'b00;
defparam dpb_inst_46.WRITE_MODE1 = 2'b00;
defparam dpb_inst_46.BIT_WIDTH_0 = 2;
defparam dpb_inst_46.BIT_WIDTH_1 = 2;
defparam dpb_inst_46.BLK_SEL_0 = 3'b010;
defparam dpb_inst_46.BLK_SEL_1 = 3'b010;
defparam dpb_inst_46.RESET_MODE = "SYNC";

DPB dpb_inst_47 (
    .DOA({dpb_inst_47_douta_w[13:0],dpb_inst_47_douta[30:29]}),
    .DOB({dpb_inst_47_doutb_w[13:0],dpb_inst_47_doutb[30:29]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[30:29]}),
    .ADB({adb[12:0],gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[30:29]})
);

defparam dpb_inst_47.READ_MODE0 = 1'b0;
defparam dpb_inst_47.READ_MODE1 = 1'b0;
defparam dpb_inst_47.WRITE_MODE0 = 2'b00;
defparam dpb_inst_47.WRITE_MODE1 = 2'b00;
defparam dpb_inst_47.BIT_WIDTH_0 = 2;
defparam dpb_inst_47.BIT_WIDTH_1 = 2;
defparam dpb_inst_47.BLK_SEL_0 = 3'b010;
defparam dpb_inst_47.BLK_SEL_1 = 3'b010;
defparam dpb_inst_47.RESET_MODE = "SYNC";

DPB dpb_inst_48 (
    .DOA({dpb_inst_48_douta_w[11:0],dpb_inst_48_douta[30:27]}),
    .DOB({dpb_inst_48_doutb_w[11:0],dpb_inst_48_doutb[30:27]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[30:27]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[30:27]})
);

defparam dpb_inst_48.READ_MODE0 = 1'b0;
defparam dpb_inst_48.READ_MODE1 = 1'b0;
defparam dpb_inst_48.WRITE_MODE0 = 2'b00;
defparam dpb_inst_48.WRITE_MODE1 = 2'b00;
defparam dpb_inst_48.BIT_WIDTH_0 = 4;
defparam dpb_inst_48.BIT_WIDTH_1 = 4;
defparam dpb_inst_48.BLK_SEL_0 = 3'b110;
defparam dpb_inst_48.BLK_SEL_1 = 3'b110;
defparam dpb_inst_48.RESET_MODE = "SYNC";

DPB dpb_inst_49 (
    .DOA({dpb_inst_49_douta_w[14:0],dpb_inst_49_douta[31]}),
    .DOB({dpb_inst_49_doutb_w[14:0],dpb_inst_49_doutb[31]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[31]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[31]})
);

defparam dpb_inst_49.READ_MODE0 = 1'b0;
defparam dpb_inst_49.READ_MODE1 = 1'b0;
defparam dpb_inst_49.WRITE_MODE0 = 2'b00;
defparam dpb_inst_49.WRITE_MODE1 = 2'b00;
defparam dpb_inst_49.BIT_WIDTH_0 = 1;
defparam dpb_inst_49.BIT_WIDTH_1 = 1;
defparam dpb_inst_49.BLK_SEL_0 = 3'b000;
defparam dpb_inst_49.BLK_SEL_1 = 3'b000;
defparam dpb_inst_49.RESET_MODE = "SYNC";

DPB dpb_inst_50 (
    .DOA({dpb_inst_50_douta_w[14:0],dpb_inst_50_douta[31]}),
    .DOB({dpb_inst_50_doutb_w[14:0],dpb_inst_50_doutb[31]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[31]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[31]})
);

defparam dpb_inst_50.READ_MODE0 = 1'b0;
defparam dpb_inst_50.READ_MODE1 = 1'b0;
defparam dpb_inst_50.WRITE_MODE0 = 2'b00;
defparam dpb_inst_50.WRITE_MODE1 = 2'b00;
defparam dpb_inst_50.BIT_WIDTH_0 = 1;
defparam dpb_inst_50.BIT_WIDTH_1 = 1;
defparam dpb_inst_50.BLK_SEL_0 = 3'b001;
defparam dpb_inst_50.BLK_SEL_1 = 3'b001;
defparam dpb_inst_50.RESET_MODE = "SYNC";

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(ada[14]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_1 (
  .Q(dff_q_1),
  .D(ada[13]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_2 (
  .Q(dff_q_2),
  .D(ada[12]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_3 (
  .Q(dff_q_3),
  .D(ada[11]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_4 (
  .Q(dff_q_4),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_5 (
  .Q(dff_q_5),
  .D(adb[13]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_6 (
  .Q(dff_q_6),
  .D(adb[12]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_7 (
  .Q(dff_q_7),
  .D(adb[11]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(dpx9b_inst_0_douta[0]),
  .I1(dpx9b_inst_1_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(dpx9b_inst_2_douta[0]),
  .I1(dpx9b_inst_3_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(dpx9b_inst_4_douta[0]),
  .I1(dpx9b_inst_5_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(dpx9b_inst_6_douta[0]),
  .I1(dpx9b_inst_7_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(dpx9b_inst_8_douta[0]),
  .I1(dpx9b_inst_9_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(dpx9b_inst_10_douta[0]),
  .I1(dpx9b_inst_11_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(dpx9b_inst_12_douta[0]),
  .I1(dpx9b_inst_13_douta[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_2)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_2)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_2)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(mux_o_7),
  .I1(mux_o_8),
  .S0(dff_q_1)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_9),
  .I1(mux_o_6),
  .S0(dff_q_1)
);
MUX2 mux_inst_13 (
  .O(douta[0]),
  .I0(mux_o_11),
  .I1(mux_o_12),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(dpx9b_inst_0_douta[1]),
  .I1(dpx9b_inst_1_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(dpx9b_inst_2_douta[1]),
  .I1(dpx9b_inst_3_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(dpx9b_inst_4_douta[1]),
  .I1(dpx9b_inst_5_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(dpx9b_inst_6_douta[1]),
  .I1(dpx9b_inst_7_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(dpx9b_inst_8_douta[1]),
  .I1(dpx9b_inst_9_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(dpx9b_inst_10_douta[1]),
  .I1(dpx9b_inst_11_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(dpx9b_inst_12_douta[1]),
  .I1(dpx9b_inst_13_douta[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(dff_q_2)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_2)
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(dff_q_2)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(dff_q_1)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_23),
  .I1(mux_o_20),
  .S0(dff_q_1)
);
MUX2 mux_inst_27 (
  .O(douta[1]),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(dff_q_0)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(dpx9b_inst_0_douta[2]),
  .I1(dpx9b_inst_1_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(dpx9b_inst_2_douta[2]),
  .I1(dpx9b_inst_3_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(dpx9b_inst_4_douta[2]),
  .I1(dpx9b_inst_5_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(dpx9b_inst_6_douta[2]),
  .I1(dpx9b_inst_7_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(dpx9b_inst_8_douta[2]),
  .I1(dpx9b_inst_9_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(dpx9b_inst_10_douta[2]),
  .I1(dpx9b_inst_11_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(dpx9b_inst_12_douta[2]),
  .I1(dpx9b_inst_13_douta[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(dff_q_2)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(dff_q_2)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(dff_q_2)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(dff_q_1)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_37),
  .I1(mux_o_34),
  .S0(dff_q_1)
);
MUX2 mux_inst_41 (
  .O(douta[2]),
  .I0(mux_o_39),
  .I1(mux_o_40),
  .S0(dff_q_0)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(dpx9b_inst_0_douta[3]),
  .I1(dpx9b_inst_1_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(dpx9b_inst_2_douta[3]),
  .I1(dpx9b_inst_3_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(dpx9b_inst_4_douta[3]),
  .I1(dpx9b_inst_5_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(dpx9b_inst_6_douta[3]),
  .I1(dpx9b_inst_7_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(dpx9b_inst_8_douta[3]),
  .I1(dpx9b_inst_9_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(dpx9b_inst_10_douta[3]),
  .I1(dpx9b_inst_11_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(dpx9b_inst_12_douta[3]),
  .I1(dpx9b_inst_13_douta[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(dff_q_2)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(mux_o_44),
  .I1(mux_o_45),
  .S0(dff_q_2)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(mux_o_46),
  .I1(mux_o_47),
  .S0(dff_q_2)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(dff_q_1)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_51),
  .I1(mux_o_48),
  .S0(dff_q_1)
);
MUX2 mux_inst_55 (
  .O(douta[3]),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(dff_q_0)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(dpx9b_inst_0_douta[4]),
  .I1(dpx9b_inst_1_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(dpx9b_inst_2_douta[4]),
  .I1(dpx9b_inst_3_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(dpx9b_inst_4_douta[4]),
  .I1(dpx9b_inst_5_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(dpx9b_inst_6_douta[4]),
  .I1(dpx9b_inst_7_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(dpx9b_inst_8_douta[4]),
  .I1(dpx9b_inst_9_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(dpx9b_inst_10_douta[4]),
  .I1(dpx9b_inst_11_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(dpx9b_inst_12_douta[4]),
  .I1(dpx9b_inst_13_douta[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(mux_o_56),
  .I1(mux_o_57),
  .S0(dff_q_2)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(mux_o_58),
  .I1(mux_o_59),
  .S0(dff_q_2)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(dff_q_2)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(mux_o_63),
  .I1(mux_o_64),
  .S0(dff_q_1)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(mux_o_65),
  .I1(mux_o_62),
  .S0(dff_q_1)
);
MUX2 mux_inst_69 (
  .O(douta[4]),
  .I0(mux_o_67),
  .I1(mux_o_68),
  .S0(dff_q_0)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(dpx9b_inst_0_douta[5]),
  .I1(dpx9b_inst_1_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(dpx9b_inst_2_douta[5]),
  .I1(dpx9b_inst_3_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(dpx9b_inst_4_douta[5]),
  .I1(dpx9b_inst_5_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(dpx9b_inst_6_douta[5]),
  .I1(dpx9b_inst_7_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(dpx9b_inst_8_douta[5]),
  .I1(dpx9b_inst_9_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(dpx9b_inst_10_douta[5]),
  .I1(dpx9b_inst_11_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(dpx9b_inst_12_douta[5]),
  .I1(dpx9b_inst_13_douta[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_2)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(dff_q_2)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(mux_o_74),
  .I1(mux_o_75),
  .S0(dff_q_2)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(dff_q_1)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(mux_o_79),
  .I1(mux_o_76),
  .S0(dff_q_1)
);
MUX2 mux_inst_83 (
  .O(douta[5]),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_0)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(dpx9b_inst_0_douta[6]),
  .I1(dpx9b_inst_1_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(dpx9b_inst_2_douta[6]),
  .I1(dpx9b_inst_3_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(dpx9b_inst_4_douta[6]),
  .I1(dpx9b_inst_5_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(dpx9b_inst_6_douta[6]),
  .I1(dpx9b_inst_7_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(dpx9b_inst_8_douta[6]),
  .I1(dpx9b_inst_9_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(dpx9b_inst_10_douta[6]),
  .I1(dpx9b_inst_11_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(dpx9b_inst_12_douta[6]),
  .I1(dpx9b_inst_13_douta[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_84),
  .I1(mux_o_85),
  .S0(dff_q_2)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(mux_o_86),
  .I1(mux_o_87),
  .S0(dff_q_2)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(dff_q_2)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_91),
  .I1(mux_o_92),
  .S0(dff_q_1)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(mux_o_93),
  .I1(mux_o_90),
  .S0(dff_q_1)
);
MUX2 mux_inst_97 (
  .O(douta[6]),
  .I0(mux_o_95),
  .I1(mux_o_96),
  .S0(dff_q_0)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(dpx9b_inst_0_douta[7]),
  .I1(dpx9b_inst_1_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(dpx9b_inst_2_douta[7]),
  .I1(dpx9b_inst_3_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(dpx9b_inst_4_douta[7]),
  .I1(dpx9b_inst_5_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(dpx9b_inst_6_douta[7]),
  .I1(dpx9b_inst_7_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(dpx9b_inst_8_douta[7]),
  .I1(dpx9b_inst_9_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(dpx9b_inst_10_douta[7]),
  .I1(dpx9b_inst_11_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(dpx9b_inst_12_douta[7]),
  .I1(dpx9b_inst_13_douta[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(dff_q_2)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(dff_q_2)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(dff_q_2)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(dff_q_1)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_107),
  .I1(mux_o_104),
  .S0(dff_q_1)
);
MUX2 mux_inst_111 (
  .O(douta[7]),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(dff_q_0)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(dpx9b_inst_0_douta[8]),
  .I1(dpx9b_inst_1_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(dpx9b_inst_2_douta[8]),
  .I1(dpx9b_inst_3_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(dpx9b_inst_4_douta[8]),
  .I1(dpx9b_inst_5_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(dpx9b_inst_6_douta[8]),
  .I1(dpx9b_inst_7_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(dpx9b_inst_8_douta[8]),
  .I1(dpx9b_inst_9_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(dpx9b_inst_10_douta[8]),
  .I1(dpx9b_inst_11_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(dpx9b_inst_12_douta[8]),
  .I1(dpx9b_inst_13_douta[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(mux_o_112),
  .I1(mux_o_113),
  .S0(dff_q_2)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(mux_o_114),
  .I1(mux_o_115),
  .S0(dff_q_2)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(mux_o_116),
  .I1(mux_o_117),
  .S0(dff_q_2)
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(mux_o_119),
  .I1(mux_o_120),
  .S0(dff_q_1)
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(mux_o_121),
  .I1(mux_o_118),
  .S0(dff_q_1)
);
MUX2 mux_inst_125 (
  .O(douta[8]),
  .I0(mux_o_123),
  .I1(mux_o_124),
  .S0(dff_q_0)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(dpx9b_inst_14_douta[9]),
  .I1(dpx9b_inst_15_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(dpx9b_inst_16_douta[9]),
  .I1(dpx9b_inst_17_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(dpx9b_inst_18_douta[9]),
  .I1(dpx9b_inst_19_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(dpx9b_inst_20_douta[9]),
  .I1(dpx9b_inst_21_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(dpx9b_inst_22_douta[9]),
  .I1(dpx9b_inst_23_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(dpx9b_inst_24_douta[9]),
  .I1(dpx9b_inst_25_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(dpx9b_inst_26_douta[9]),
  .I1(dpx9b_inst_27_douta[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(dff_q_2)
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(dff_q_2)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_2)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(mux_o_133),
  .I1(mux_o_134),
  .S0(dff_q_1)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(mux_o_135),
  .I1(mux_o_132),
  .S0(dff_q_1)
);
MUX2 mux_inst_139 (
  .O(douta[9]),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(dff_q_0)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(dpx9b_inst_14_douta[10]),
  .I1(dpx9b_inst_15_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(dpx9b_inst_16_douta[10]),
  .I1(dpx9b_inst_17_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(dpx9b_inst_18_douta[10]),
  .I1(dpx9b_inst_19_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(dpx9b_inst_20_douta[10]),
  .I1(dpx9b_inst_21_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(dpx9b_inst_22_douta[10]),
  .I1(dpx9b_inst_23_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(dpx9b_inst_24_douta[10]),
  .I1(dpx9b_inst_25_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(dpx9b_inst_26_douta[10]),
  .I1(dpx9b_inst_27_douta[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_140),
  .I1(mux_o_141),
  .S0(dff_q_2)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(dff_q_2)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(dff_q_2)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(mux_o_147),
  .I1(mux_o_148),
  .S0(dff_q_1)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(mux_o_149),
  .I1(mux_o_146),
  .S0(dff_q_1)
);
MUX2 mux_inst_153 (
  .O(douta[10]),
  .I0(mux_o_151),
  .I1(mux_o_152),
  .S0(dff_q_0)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(dpx9b_inst_14_douta[11]),
  .I1(dpx9b_inst_15_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(dpx9b_inst_16_douta[11]),
  .I1(dpx9b_inst_17_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(dpx9b_inst_18_douta[11]),
  .I1(dpx9b_inst_19_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(dpx9b_inst_20_douta[11]),
  .I1(dpx9b_inst_21_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(dpx9b_inst_22_douta[11]),
  .I1(dpx9b_inst_23_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(dpx9b_inst_24_douta[11]),
  .I1(dpx9b_inst_25_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(dpx9b_inst_26_douta[11]),
  .I1(dpx9b_inst_27_douta[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(dff_q_2)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(dff_q_2)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(dff_q_2)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(mux_o_161),
  .I1(mux_o_162),
  .S0(dff_q_1)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(mux_o_163),
  .I1(mux_o_160),
  .S0(dff_q_1)
);
MUX2 mux_inst_167 (
  .O(douta[11]),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(dff_q_0)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(dpx9b_inst_14_douta[12]),
  .I1(dpx9b_inst_15_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(dpx9b_inst_16_douta[12]),
  .I1(dpx9b_inst_17_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(dpx9b_inst_18_douta[12]),
  .I1(dpx9b_inst_19_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(dpx9b_inst_20_douta[12]),
  .I1(dpx9b_inst_21_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(dpx9b_inst_22_douta[12]),
  .I1(dpx9b_inst_23_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(dpx9b_inst_24_douta[12]),
  .I1(dpx9b_inst_25_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(dpx9b_inst_26_douta[12]),
  .I1(dpx9b_inst_27_douta[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(mux_o_168),
  .I1(mux_o_169),
  .S0(dff_q_2)
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(mux_o_170),
  .I1(mux_o_171),
  .S0(dff_q_2)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_172),
  .I1(mux_o_173),
  .S0(dff_q_2)
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(dff_q_1)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(mux_o_177),
  .I1(mux_o_174),
  .S0(dff_q_1)
);
MUX2 mux_inst_181 (
  .O(douta[12]),
  .I0(mux_o_179),
  .I1(mux_o_180),
  .S0(dff_q_0)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(dpx9b_inst_14_douta[13]),
  .I1(dpx9b_inst_15_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(dpx9b_inst_16_douta[13]),
  .I1(dpx9b_inst_17_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(dpx9b_inst_18_douta[13]),
  .I1(dpx9b_inst_19_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(dpx9b_inst_20_douta[13]),
  .I1(dpx9b_inst_21_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(dpx9b_inst_22_douta[13]),
  .I1(dpx9b_inst_23_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(dpx9b_inst_24_douta[13]),
  .I1(dpx9b_inst_25_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(dpx9b_inst_26_douta[13]),
  .I1(dpx9b_inst_27_douta[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(dff_q_2)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(dff_q_2)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(dff_q_2)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(dff_q_1)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(mux_o_191),
  .I1(mux_o_188),
  .S0(dff_q_1)
);
MUX2 mux_inst_195 (
  .O(douta[13]),
  .I0(mux_o_193),
  .I1(mux_o_194),
  .S0(dff_q_0)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(dpx9b_inst_14_douta[14]),
  .I1(dpx9b_inst_15_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(dpx9b_inst_16_douta[14]),
  .I1(dpx9b_inst_17_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(dpx9b_inst_18_douta[14]),
  .I1(dpx9b_inst_19_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(dpx9b_inst_20_douta[14]),
  .I1(dpx9b_inst_21_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(dpx9b_inst_22_douta[14]),
  .I1(dpx9b_inst_23_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(dpx9b_inst_24_douta[14]),
  .I1(dpx9b_inst_25_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(dpx9b_inst_26_douta[14]),
  .I1(dpx9b_inst_27_douta[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(dff_q_2)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(dff_q_2)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_200),
  .I1(mux_o_201),
  .S0(dff_q_2)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(dff_q_1)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_205),
  .I1(mux_o_202),
  .S0(dff_q_1)
);
MUX2 mux_inst_209 (
  .O(douta[14]),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(dff_q_0)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(dpx9b_inst_14_douta[15]),
  .I1(dpx9b_inst_15_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(dpx9b_inst_16_douta[15]),
  .I1(dpx9b_inst_17_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(dpx9b_inst_18_douta[15]),
  .I1(dpx9b_inst_19_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(dpx9b_inst_20_douta[15]),
  .I1(dpx9b_inst_21_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(dpx9b_inst_22_douta[15]),
  .I1(dpx9b_inst_23_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(dpx9b_inst_24_douta[15]),
  .I1(dpx9b_inst_25_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(dpx9b_inst_26_douta[15]),
  .I1(dpx9b_inst_27_douta[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(dff_q_2)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(dff_q_2)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(dff_q_2)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(dff_q_1)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_219),
  .I1(mux_o_216),
  .S0(dff_q_1)
);
MUX2 mux_inst_223 (
  .O(douta[15]),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(dff_q_0)
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(dpx9b_inst_14_douta[16]),
  .I1(dpx9b_inst_15_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(dpx9b_inst_16_douta[16]),
  .I1(dpx9b_inst_17_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(dpx9b_inst_18_douta[16]),
  .I1(dpx9b_inst_19_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(dpx9b_inst_20_douta[16]),
  .I1(dpx9b_inst_21_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(dpx9b_inst_22_douta[16]),
  .I1(dpx9b_inst_23_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(dpx9b_inst_24_douta[16]),
  .I1(dpx9b_inst_25_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(dpx9b_inst_26_douta[16]),
  .I1(dpx9b_inst_27_douta[16]),
  .S0(dff_q_3)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(mux_o_224),
  .I1(mux_o_225),
  .S0(dff_q_2)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(mux_o_226),
  .I1(mux_o_227),
  .S0(dff_q_2)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_228),
  .I1(mux_o_229),
  .S0(dff_q_2)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_1)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_233),
  .I1(mux_o_230),
  .S0(dff_q_1)
);
MUX2 mux_inst_237 (
  .O(douta[16]),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_0)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(dpx9b_inst_14_douta[17]),
  .I1(dpx9b_inst_15_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(dpx9b_inst_16_douta[17]),
  .I1(dpx9b_inst_17_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(dpx9b_inst_18_douta[17]),
  .I1(dpx9b_inst_19_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(dpx9b_inst_20_douta[17]),
  .I1(dpx9b_inst_21_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(dpx9b_inst_22_douta[17]),
  .I1(dpx9b_inst_23_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(dpx9b_inst_24_douta[17]),
  .I1(dpx9b_inst_25_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(dpx9b_inst_26_douta[17]),
  .I1(dpx9b_inst_27_douta[17]),
  .S0(dff_q_3)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(mux_o_238),
  .I1(mux_o_239),
  .S0(dff_q_2)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_240),
  .I1(mux_o_241),
  .S0(dff_q_2)
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(mux_o_242),
  .I1(mux_o_243),
  .S0(dff_q_2)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_245),
  .I1(mux_o_246),
  .S0(dff_q_1)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_247),
  .I1(mux_o_244),
  .S0(dff_q_1)
);
MUX2 mux_inst_251 (
  .O(douta[17]),
  .I0(mux_o_249),
  .I1(mux_o_250),
  .S0(dff_q_0)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(dpx9b_inst_28_douta[18]),
  .I1(dpx9b_inst_29_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(dpx9b_inst_30_douta[18]),
  .I1(dpx9b_inst_31_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(dpx9b_inst_32_douta[18]),
  .I1(dpx9b_inst_33_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(dpx9b_inst_34_douta[18]),
  .I1(dpx9b_inst_35_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(dpx9b_inst_36_douta[18]),
  .I1(dpx9b_inst_37_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(dpx9b_inst_38_douta[18]),
  .I1(dpx9b_inst_39_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(dpx9b_inst_40_douta[18]),
  .I1(dpx9b_inst_41_douta[18]),
  .S0(dff_q_3)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(dff_q_2)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(mux_o_254),
  .I1(mux_o_255),
  .S0(dff_q_2)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(mux_o_256),
  .I1(mux_o_257),
  .S0(dff_q_2)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(mux_o_259),
  .I1(mux_o_260),
  .S0(dff_q_1)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(mux_o_261),
  .I1(mux_o_258),
  .S0(dff_q_1)
);
MUX2 mux_inst_265 (
  .O(douta[18]),
  .I0(mux_o_263),
  .I1(mux_o_264),
  .S0(dff_q_0)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(dpx9b_inst_28_douta[19]),
  .I1(dpx9b_inst_29_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(dpx9b_inst_30_douta[19]),
  .I1(dpx9b_inst_31_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(dpx9b_inst_32_douta[19]),
  .I1(dpx9b_inst_33_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(dpx9b_inst_34_douta[19]),
  .I1(dpx9b_inst_35_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(dpx9b_inst_36_douta[19]),
  .I1(dpx9b_inst_37_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(dpx9b_inst_38_douta[19]),
  .I1(dpx9b_inst_39_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(dpx9b_inst_40_douta[19]),
  .I1(dpx9b_inst_41_douta[19]),
  .S0(dff_q_3)
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(dff_q_2)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(dff_q_2)
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(dff_q_2)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(mux_o_273),
  .I1(mux_o_274),
  .S0(dff_q_1)
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(mux_o_275),
  .I1(mux_o_272),
  .S0(dff_q_1)
);
MUX2 mux_inst_279 (
  .O(douta[19]),
  .I0(mux_o_277),
  .I1(mux_o_278),
  .S0(dff_q_0)
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(dpx9b_inst_28_douta[20]),
  .I1(dpx9b_inst_29_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(dpx9b_inst_30_douta[20]),
  .I1(dpx9b_inst_31_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(dpx9b_inst_32_douta[20]),
  .I1(dpx9b_inst_33_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(dpx9b_inst_34_douta[20]),
  .I1(dpx9b_inst_35_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(dpx9b_inst_36_douta[20]),
  .I1(dpx9b_inst_37_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(dpx9b_inst_38_douta[20]),
  .I1(dpx9b_inst_39_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(dpx9b_inst_40_douta[20]),
  .I1(dpx9b_inst_41_douta[20]),
  .S0(dff_q_3)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(dff_q_2)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(dff_q_2)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(mux_o_284),
  .I1(mux_o_285),
  .S0(dff_q_2)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(dff_q_1)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(mux_o_289),
  .I1(mux_o_286),
  .S0(dff_q_1)
);
MUX2 mux_inst_293 (
  .O(douta[20]),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(dff_q_0)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(dpx9b_inst_28_douta[21]),
  .I1(dpx9b_inst_29_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(dpx9b_inst_30_douta[21]),
  .I1(dpx9b_inst_31_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(dpx9b_inst_32_douta[21]),
  .I1(dpx9b_inst_33_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(dpx9b_inst_34_douta[21]),
  .I1(dpx9b_inst_35_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(dpx9b_inst_36_douta[21]),
  .I1(dpx9b_inst_37_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(dpx9b_inst_38_douta[21]),
  .I1(dpx9b_inst_39_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(dpx9b_inst_40_douta[21]),
  .I1(dpx9b_inst_41_douta[21]),
  .S0(dff_q_3)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(mux_o_294),
  .I1(mux_o_295),
  .S0(dff_q_2)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(mux_o_296),
  .I1(mux_o_297),
  .S0(dff_q_2)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(dff_q_2)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(mux_o_301),
  .I1(mux_o_302),
  .S0(dff_q_1)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(mux_o_303),
  .I1(mux_o_300),
  .S0(dff_q_1)
);
MUX2 mux_inst_307 (
  .O(douta[21]),
  .I0(mux_o_305),
  .I1(mux_o_306),
  .S0(dff_q_0)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(dpx9b_inst_28_douta[22]),
  .I1(dpx9b_inst_29_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(dpx9b_inst_30_douta[22]),
  .I1(dpx9b_inst_31_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(dpx9b_inst_32_douta[22]),
  .I1(dpx9b_inst_33_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(dpx9b_inst_34_douta[22]),
  .I1(dpx9b_inst_35_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(dpx9b_inst_36_douta[22]),
  .I1(dpx9b_inst_37_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(dpx9b_inst_38_douta[22]),
  .I1(dpx9b_inst_39_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_314 (
  .O(mux_o_314),
  .I0(dpx9b_inst_40_douta[22]),
  .I1(dpx9b_inst_41_douta[22]),
  .S0(dff_q_3)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(dff_q_2)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(dff_q_2)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(dff_q_2)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(mux_o_315),
  .I1(mux_o_316),
  .S0(dff_q_1)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(mux_o_317),
  .I1(mux_o_314),
  .S0(dff_q_1)
);
MUX2 mux_inst_321 (
  .O(douta[22]),
  .I0(mux_o_319),
  .I1(mux_o_320),
  .S0(dff_q_0)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(dpx9b_inst_28_douta[23]),
  .I1(dpx9b_inst_29_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(dpx9b_inst_30_douta[23]),
  .I1(dpx9b_inst_31_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(dpx9b_inst_32_douta[23]),
  .I1(dpx9b_inst_33_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(dpx9b_inst_34_douta[23]),
  .I1(dpx9b_inst_35_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(dpx9b_inst_36_douta[23]),
  .I1(dpx9b_inst_37_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(dpx9b_inst_38_douta[23]),
  .I1(dpx9b_inst_39_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(dpx9b_inst_40_douta[23]),
  .I1(dpx9b_inst_41_douta[23]),
  .S0(dff_q_3)
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(mux_o_322),
  .I1(mux_o_323),
  .S0(dff_q_2)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(mux_o_324),
  .I1(mux_o_325),
  .S0(dff_q_2)
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(mux_o_326),
  .I1(mux_o_327),
  .S0(dff_q_2)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(mux_o_329),
  .I1(mux_o_330),
  .S0(dff_q_1)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(mux_o_331),
  .I1(mux_o_328),
  .S0(dff_q_1)
);
MUX2 mux_inst_335 (
  .O(douta[23]),
  .I0(mux_o_333),
  .I1(mux_o_334),
  .S0(dff_q_0)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(dpx9b_inst_28_douta[24]),
  .I1(dpx9b_inst_29_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(dpx9b_inst_30_douta[24]),
  .I1(dpx9b_inst_31_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(dpx9b_inst_32_douta[24]),
  .I1(dpx9b_inst_33_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(dpx9b_inst_34_douta[24]),
  .I1(dpx9b_inst_35_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(dpx9b_inst_36_douta[24]),
  .I1(dpx9b_inst_37_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(dpx9b_inst_38_douta[24]),
  .I1(dpx9b_inst_39_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(dpx9b_inst_40_douta[24]),
  .I1(dpx9b_inst_41_douta[24]),
  .S0(dff_q_3)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(dff_q_2)
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(dff_q_2)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(mux_o_340),
  .I1(mux_o_341),
  .S0(dff_q_2)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(mux_o_343),
  .I1(mux_o_344),
  .S0(dff_q_1)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(mux_o_345),
  .I1(mux_o_342),
  .S0(dff_q_1)
);
MUX2 mux_inst_349 (
  .O(douta[24]),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_0)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(dpx9b_inst_28_douta[25]),
  .I1(dpx9b_inst_29_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(dpx9b_inst_30_douta[25]),
  .I1(dpx9b_inst_31_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(dpx9b_inst_32_douta[25]),
  .I1(dpx9b_inst_33_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(dpx9b_inst_34_douta[25]),
  .I1(dpx9b_inst_35_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(dpx9b_inst_36_douta[25]),
  .I1(dpx9b_inst_37_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(dpx9b_inst_38_douta[25]),
  .I1(dpx9b_inst_39_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(dpx9b_inst_40_douta[25]),
  .I1(dpx9b_inst_41_douta[25]),
  .S0(dff_q_3)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_350),
  .I1(mux_o_351),
  .S0(dff_q_2)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_352),
  .I1(mux_o_353),
  .S0(dff_q_2)
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_354),
  .I1(mux_o_355),
  .S0(dff_q_2)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_1)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_359),
  .I1(mux_o_356),
  .S0(dff_q_1)
);
MUX2 mux_inst_363 (
  .O(douta[25]),
  .I0(mux_o_361),
  .I1(mux_o_362),
  .S0(dff_q_0)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(dpx9b_inst_28_douta[26]),
  .I1(dpx9b_inst_29_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(dpx9b_inst_30_douta[26]),
  .I1(dpx9b_inst_31_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(dpx9b_inst_32_douta[26]),
  .I1(dpx9b_inst_33_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(dpx9b_inst_34_douta[26]),
  .I1(dpx9b_inst_35_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(dpx9b_inst_36_douta[26]),
  .I1(dpx9b_inst_37_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(dpx9b_inst_38_douta[26]),
  .I1(dpx9b_inst_39_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(dpx9b_inst_40_douta[26]),
  .I1(dpx9b_inst_41_douta[26]),
  .S0(dff_q_3)
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(mux_o_364),
  .I1(mux_o_365),
  .S0(dff_q_2)
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(mux_o_366),
  .I1(mux_o_367),
  .S0(dff_q_2)
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(mux_o_368),
  .I1(mux_o_369),
  .S0(dff_q_2)
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(mux_o_371),
  .I1(mux_o_372),
  .S0(dff_q_1)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(mux_o_373),
  .I1(mux_o_370),
  .S0(dff_q_1)
);
MUX2 mux_inst_377 (
  .O(douta[26]),
  .I0(mux_o_375),
  .I1(mux_o_376),
  .S0(dff_q_0)
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(dpb_inst_46_douta[27]),
  .I1(dpb_inst_48_douta[27]),
  .S0(dff_q_1)
);
MUX2 mux_inst_386 (
  .O(douta[27]),
  .I0(dpb_inst_42_douta[27]),
  .I1(mux_o_385),
  .S0(dff_q_0)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(dpb_inst_46_douta[28]),
  .I1(dpb_inst_48_douta[28]),
  .S0(dff_q_1)
);
MUX2 mux_inst_395 (
  .O(douta[28]),
  .I0(dpb_inst_43_douta[28]),
  .I1(mux_o_394),
  .S0(dff_q_0)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(dpb_inst_47_douta[29]),
  .I1(dpb_inst_48_douta[29]),
  .S0(dff_q_1)
);
MUX2 mux_inst_404 (
  .O(douta[29]),
  .I0(dpb_inst_44_douta[29]),
  .I1(mux_o_403),
  .S0(dff_q_0)
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(dpb_inst_47_douta[30]),
  .I1(dpb_inst_48_douta[30]),
  .S0(dff_q_1)
);
MUX2 mux_inst_413 (
  .O(douta[30]),
  .I0(dpb_inst_45_douta[30]),
  .I1(mux_o_412),
  .S0(dff_q_0)
);
MUX2 mux_inst_420 (
  .O(douta[31]),
  .I0(dpb_inst_49_douta[31]),
  .I1(dpb_inst_50_douta[31]),
  .S0(dff_q_0)
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(dpx9b_inst_0_doutb[0]),
  .I1(dpx9b_inst_1_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(dpx9b_inst_2_doutb[0]),
  .I1(dpx9b_inst_3_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(dpx9b_inst_4_doutb[0]),
  .I1(dpx9b_inst_5_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(dpx9b_inst_6_doutb[0]),
  .I1(dpx9b_inst_7_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(dpx9b_inst_8_doutb[0]),
  .I1(dpx9b_inst_9_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(dpx9b_inst_10_doutb[0]),
  .I1(dpx9b_inst_11_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(dpx9b_inst_12_doutb[0]),
  .I1(dpx9b_inst_13_doutb[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(mux_o_421),
  .I1(mux_o_422),
  .S0(dff_q_6)
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(mux_o_423),
  .I1(mux_o_424),
  .S0(dff_q_6)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(mux_o_425),
  .I1(mux_o_426),
  .S0(dff_q_6)
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(mux_o_428),
  .I1(mux_o_429),
  .S0(dff_q_5)
);
MUX2 mux_inst_433 (
  .O(mux_o_433),
  .I0(mux_o_430),
  .I1(mux_o_427),
  .S0(dff_q_5)
);
MUX2 mux_inst_434 (
  .O(doutb[0]),
  .I0(mux_o_432),
  .I1(mux_o_433),
  .S0(dff_q_4)
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(dpx9b_inst_0_doutb[1]),
  .I1(dpx9b_inst_1_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(dpx9b_inst_2_doutb[1]),
  .I1(dpx9b_inst_3_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(dpx9b_inst_4_doutb[1]),
  .I1(dpx9b_inst_5_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(dpx9b_inst_6_doutb[1]),
  .I1(dpx9b_inst_7_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(dpx9b_inst_8_doutb[1]),
  .I1(dpx9b_inst_9_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(dpx9b_inst_10_doutb[1]),
  .I1(dpx9b_inst_11_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(dpx9b_inst_12_doutb[1]),
  .I1(dpx9b_inst_13_doutb[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(mux_o_435),
  .I1(mux_o_436),
  .S0(dff_q_6)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(mux_o_437),
  .I1(mux_o_438),
  .S0(dff_q_6)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(mux_o_439),
  .I1(mux_o_440),
  .S0(dff_q_6)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(mux_o_442),
  .I1(mux_o_443),
  .S0(dff_q_5)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(mux_o_444),
  .I1(mux_o_441),
  .S0(dff_q_5)
);
MUX2 mux_inst_448 (
  .O(doutb[1]),
  .I0(mux_o_446),
  .I1(mux_o_447),
  .S0(dff_q_4)
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(dpx9b_inst_0_doutb[2]),
  .I1(dpx9b_inst_1_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(dpx9b_inst_2_doutb[2]),
  .I1(dpx9b_inst_3_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(dpx9b_inst_4_doutb[2]),
  .I1(dpx9b_inst_5_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(dpx9b_inst_6_doutb[2]),
  .I1(dpx9b_inst_7_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(dpx9b_inst_8_doutb[2]),
  .I1(dpx9b_inst_9_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(dpx9b_inst_10_doutb[2]),
  .I1(dpx9b_inst_11_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(dpx9b_inst_12_doutb[2]),
  .I1(dpx9b_inst_13_doutb[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(mux_o_449),
  .I1(mux_o_450),
  .S0(dff_q_6)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(mux_o_451),
  .I1(mux_o_452),
  .S0(dff_q_6)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_453),
  .I1(mux_o_454),
  .S0(dff_q_6)
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(mux_o_456),
  .I1(mux_o_457),
  .S0(dff_q_5)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_458),
  .I1(mux_o_455),
  .S0(dff_q_5)
);
MUX2 mux_inst_462 (
  .O(doutb[2]),
  .I0(mux_o_460),
  .I1(mux_o_461),
  .S0(dff_q_4)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(dpx9b_inst_0_doutb[3]),
  .I1(dpx9b_inst_1_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_464 (
  .O(mux_o_464),
  .I0(dpx9b_inst_2_doutb[3]),
  .I1(dpx9b_inst_3_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(dpx9b_inst_4_doutb[3]),
  .I1(dpx9b_inst_5_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(dpx9b_inst_6_doutb[3]),
  .I1(dpx9b_inst_7_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(dpx9b_inst_8_doutb[3]),
  .I1(dpx9b_inst_9_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(dpx9b_inst_10_doutb[3]),
  .I1(dpx9b_inst_11_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(dpx9b_inst_12_doutb[3]),
  .I1(dpx9b_inst_13_doutb[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(mux_o_463),
  .I1(mux_o_464),
  .S0(dff_q_6)
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_6)
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(mux_o_467),
  .I1(mux_o_468),
  .S0(dff_q_6)
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(mux_o_470),
  .I1(mux_o_471),
  .S0(dff_q_5)
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(mux_o_472),
  .I1(mux_o_469),
  .S0(dff_q_5)
);
MUX2 mux_inst_476 (
  .O(doutb[3]),
  .I0(mux_o_474),
  .I1(mux_o_475),
  .S0(dff_q_4)
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(dpx9b_inst_0_doutb[4]),
  .I1(dpx9b_inst_1_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(dpx9b_inst_2_doutb[4]),
  .I1(dpx9b_inst_3_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_479 (
  .O(mux_o_479),
  .I0(dpx9b_inst_4_doutb[4]),
  .I1(dpx9b_inst_5_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_480 (
  .O(mux_o_480),
  .I0(dpx9b_inst_6_doutb[4]),
  .I1(dpx9b_inst_7_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_481 (
  .O(mux_o_481),
  .I0(dpx9b_inst_8_doutb[4]),
  .I1(dpx9b_inst_9_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_482 (
  .O(mux_o_482),
  .I0(dpx9b_inst_10_doutb[4]),
  .I1(dpx9b_inst_11_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_483 (
  .O(mux_o_483),
  .I0(dpx9b_inst_12_doutb[4]),
  .I1(dpx9b_inst_13_doutb[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(dff_q_6)
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(mux_o_479),
  .I1(mux_o_480),
  .S0(dff_q_6)
);
MUX2 mux_inst_486 (
  .O(mux_o_486),
  .I0(mux_o_481),
  .I1(mux_o_482),
  .S0(dff_q_6)
);
MUX2 mux_inst_488 (
  .O(mux_o_488),
  .I0(mux_o_484),
  .I1(mux_o_485),
  .S0(dff_q_5)
);
MUX2 mux_inst_489 (
  .O(mux_o_489),
  .I0(mux_o_486),
  .I1(mux_o_483),
  .S0(dff_q_5)
);
MUX2 mux_inst_490 (
  .O(doutb[4]),
  .I0(mux_o_488),
  .I1(mux_o_489),
  .S0(dff_q_4)
);
MUX2 mux_inst_491 (
  .O(mux_o_491),
  .I0(dpx9b_inst_0_doutb[5]),
  .I1(dpx9b_inst_1_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_492 (
  .O(mux_o_492),
  .I0(dpx9b_inst_2_doutb[5]),
  .I1(dpx9b_inst_3_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_493 (
  .O(mux_o_493),
  .I0(dpx9b_inst_4_doutb[5]),
  .I1(dpx9b_inst_5_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_494 (
  .O(mux_o_494),
  .I0(dpx9b_inst_6_doutb[5]),
  .I1(dpx9b_inst_7_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_495 (
  .O(mux_o_495),
  .I0(dpx9b_inst_8_doutb[5]),
  .I1(dpx9b_inst_9_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_496 (
  .O(mux_o_496),
  .I0(dpx9b_inst_10_doutb[5]),
  .I1(dpx9b_inst_11_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_497 (
  .O(mux_o_497),
  .I0(dpx9b_inst_12_doutb[5]),
  .I1(dpx9b_inst_13_doutb[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_498 (
  .O(mux_o_498),
  .I0(mux_o_491),
  .I1(mux_o_492),
  .S0(dff_q_6)
);
MUX2 mux_inst_499 (
  .O(mux_o_499),
  .I0(mux_o_493),
  .I1(mux_o_494),
  .S0(dff_q_6)
);
MUX2 mux_inst_500 (
  .O(mux_o_500),
  .I0(mux_o_495),
  .I1(mux_o_496),
  .S0(dff_q_6)
);
MUX2 mux_inst_502 (
  .O(mux_o_502),
  .I0(mux_o_498),
  .I1(mux_o_499),
  .S0(dff_q_5)
);
MUX2 mux_inst_503 (
  .O(mux_o_503),
  .I0(mux_o_500),
  .I1(mux_o_497),
  .S0(dff_q_5)
);
MUX2 mux_inst_504 (
  .O(doutb[5]),
  .I0(mux_o_502),
  .I1(mux_o_503),
  .S0(dff_q_4)
);
MUX2 mux_inst_505 (
  .O(mux_o_505),
  .I0(dpx9b_inst_0_doutb[6]),
  .I1(dpx9b_inst_1_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_506 (
  .O(mux_o_506),
  .I0(dpx9b_inst_2_doutb[6]),
  .I1(dpx9b_inst_3_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_507 (
  .O(mux_o_507),
  .I0(dpx9b_inst_4_doutb[6]),
  .I1(dpx9b_inst_5_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_508 (
  .O(mux_o_508),
  .I0(dpx9b_inst_6_doutb[6]),
  .I1(dpx9b_inst_7_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_509 (
  .O(mux_o_509),
  .I0(dpx9b_inst_8_doutb[6]),
  .I1(dpx9b_inst_9_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_510 (
  .O(mux_o_510),
  .I0(dpx9b_inst_10_doutb[6]),
  .I1(dpx9b_inst_11_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_511 (
  .O(mux_o_511),
  .I0(dpx9b_inst_12_doutb[6]),
  .I1(dpx9b_inst_13_doutb[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_512 (
  .O(mux_o_512),
  .I0(mux_o_505),
  .I1(mux_o_506),
  .S0(dff_q_6)
);
MUX2 mux_inst_513 (
  .O(mux_o_513),
  .I0(mux_o_507),
  .I1(mux_o_508),
  .S0(dff_q_6)
);
MUX2 mux_inst_514 (
  .O(mux_o_514),
  .I0(mux_o_509),
  .I1(mux_o_510),
  .S0(dff_q_6)
);
MUX2 mux_inst_516 (
  .O(mux_o_516),
  .I0(mux_o_512),
  .I1(mux_o_513),
  .S0(dff_q_5)
);
MUX2 mux_inst_517 (
  .O(mux_o_517),
  .I0(mux_o_514),
  .I1(mux_o_511),
  .S0(dff_q_5)
);
MUX2 mux_inst_518 (
  .O(doutb[6]),
  .I0(mux_o_516),
  .I1(mux_o_517),
  .S0(dff_q_4)
);
MUX2 mux_inst_519 (
  .O(mux_o_519),
  .I0(dpx9b_inst_0_doutb[7]),
  .I1(dpx9b_inst_1_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_520 (
  .O(mux_o_520),
  .I0(dpx9b_inst_2_doutb[7]),
  .I1(dpx9b_inst_3_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_521 (
  .O(mux_o_521),
  .I0(dpx9b_inst_4_doutb[7]),
  .I1(dpx9b_inst_5_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(dpx9b_inst_6_doutb[7]),
  .I1(dpx9b_inst_7_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(dpx9b_inst_8_doutb[7]),
  .I1(dpx9b_inst_9_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_524 (
  .O(mux_o_524),
  .I0(dpx9b_inst_10_doutb[7]),
  .I1(dpx9b_inst_11_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_525 (
  .O(mux_o_525),
  .I0(dpx9b_inst_12_doutb[7]),
  .I1(dpx9b_inst_13_doutb[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_526 (
  .O(mux_o_526),
  .I0(mux_o_519),
  .I1(mux_o_520),
  .S0(dff_q_6)
);
MUX2 mux_inst_527 (
  .O(mux_o_527),
  .I0(mux_o_521),
  .I1(mux_o_522),
  .S0(dff_q_6)
);
MUX2 mux_inst_528 (
  .O(mux_o_528),
  .I0(mux_o_523),
  .I1(mux_o_524),
  .S0(dff_q_6)
);
MUX2 mux_inst_530 (
  .O(mux_o_530),
  .I0(mux_o_526),
  .I1(mux_o_527),
  .S0(dff_q_5)
);
MUX2 mux_inst_531 (
  .O(mux_o_531),
  .I0(mux_o_528),
  .I1(mux_o_525),
  .S0(dff_q_5)
);
MUX2 mux_inst_532 (
  .O(doutb[7]),
  .I0(mux_o_530),
  .I1(mux_o_531),
  .S0(dff_q_4)
);
MUX2 mux_inst_533 (
  .O(mux_o_533),
  .I0(dpx9b_inst_0_doutb[8]),
  .I1(dpx9b_inst_1_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_534 (
  .O(mux_o_534),
  .I0(dpx9b_inst_2_doutb[8]),
  .I1(dpx9b_inst_3_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_535 (
  .O(mux_o_535),
  .I0(dpx9b_inst_4_doutb[8]),
  .I1(dpx9b_inst_5_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_536 (
  .O(mux_o_536),
  .I0(dpx9b_inst_6_doutb[8]),
  .I1(dpx9b_inst_7_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_537 (
  .O(mux_o_537),
  .I0(dpx9b_inst_8_doutb[8]),
  .I1(dpx9b_inst_9_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_538 (
  .O(mux_o_538),
  .I0(dpx9b_inst_10_doutb[8]),
  .I1(dpx9b_inst_11_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_539 (
  .O(mux_o_539),
  .I0(dpx9b_inst_12_doutb[8]),
  .I1(dpx9b_inst_13_doutb[8]),
  .S0(dff_q_7)
);
MUX2 mux_inst_540 (
  .O(mux_o_540),
  .I0(mux_o_533),
  .I1(mux_o_534),
  .S0(dff_q_6)
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(mux_o_535),
  .I1(mux_o_536),
  .S0(dff_q_6)
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(mux_o_537),
  .I1(mux_o_538),
  .S0(dff_q_6)
);
MUX2 mux_inst_544 (
  .O(mux_o_544),
  .I0(mux_o_540),
  .I1(mux_o_541),
  .S0(dff_q_5)
);
MUX2 mux_inst_545 (
  .O(mux_o_545),
  .I0(mux_o_542),
  .I1(mux_o_539),
  .S0(dff_q_5)
);
MUX2 mux_inst_546 (
  .O(doutb[8]),
  .I0(mux_o_544),
  .I1(mux_o_545),
  .S0(dff_q_4)
);
MUX2 mux_inst_547 (
  .O(mux_o_547),
  .I0(dpx9b_inst_14_doutb[9]),
  .I1(dpx9b_inst_15_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_548 (
  .O(mux_o_548),
  .I0(dpx9b_inst_16_doutb[9]),
  .I1(dpx9b_inst_17_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_549 (
  .O(mux_o_549),
  .I0(dpx9b_inst_18_doutb[9]),
  .I1(dpx9b_inst_19_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_550 (
  .O(mux_o_550),
  .I0(dpx9b_inst_20_doutb[9]),
  .I1(dpx9b_inst_21_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_551 (
  .O(mux_o_551),
  .I0(dpx9b_inst_22_doutb[9]),
  .I1(dpx9b_inst_23_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_552 (
  .O(mux_o_552),
  .I0(dpx9b_inst_24_doutb[9]),
  .I1(dpx9b_inst_25_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_553 (
  .O(mux_o_553),
  .I0(dpx9b_inst_26_doutb[9]),
  .I1(dpx9b_inst_27_doutb[9]),
  .S0(dff_q_7)
);
MUX2 mux_inst_554 (
  .O(mux_o_554),
  .I0(mux_o_547),
  .I1(mux_o_548),
  .S0(dff_q_6)
);
MUX2 mux_inst_555 (
  .O(mux_o_555),
  .I0(mux_o_549),
  .I1(mux_o_550),
  .S0(dff_q_6)
);
MUX2 mux_inst_556 (
  .O(mux_o_556),
  .I0(mux_o_551),
  .I1(mux_o_552),
  .S0(dff_q_6)
);
MUX2 mux_inst_558 (
  .O(mux_o_558),
  .I0(mux_o_554),
  .I1(mux_o_555),
  .S0(dff_q_5)
);
MUX2 mux_inst_559 (
  .O(mux_o_559),
  .I0(mux_o_556),
  .I1(mux_o_553),
  .S0(dff_q_5)
);
MUX2 mux_inst_560 (
  .O(doutb[9]),
  .I0(mux_o_558),
  .I1(mux_o_559),
  .S0(dff_q_4)
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(dpx9b_inst_14_doutb[10]),
  .I1(dpx9b_inst_15_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_562 (
  .O(mux_o_562),
  .I0(dpx9b_inst_16_doutb[10]),
  .I1(dpx9b_inst_17_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_563 (
  .O(mux_o_563),
  .I0(dpx9b_inst_18_doutb[10]),
  .I1(dpx9b_inst_19_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_564 (
  .O(mux_o_564),
  .I0(dpx9b_inst_20_doutb[10]),
  .I1(dpx9b_inst_21_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_565 (
  .O(mux_o_565),
  .I0(dpx9b_inst_22_doutb[10]),
  .I1(dpx9b_inst_23_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_566 (
  .O(mux_o_566),
  .I0(dpx9b_inst_24_doutb[10]),
  .I1(dpx9b_inst_25_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_567 (
  .O(mux_o_567),
  .I0(dpx9b_inst_26_doutb[10]),
  .I1(dpx9b_inst_27_doutb[10]),
  .S0(dff_q_7)
);
MUX2 mux_inst_568 (
  .O(mux_o_568),
  .I0(mux_o_561),
  .I1(mux_o_562),
  .S0(dff_q_6)
);
MUX2 mux_inst_569 (
  .O(mux_o_569),
  .I0(mux_o_563),
  .I1(mux_o_564),
  .S0(dff_q_6)
);
MUX2 mux_inst_570 (
  .O(mux_o_570),
  .I0(mux_o_565),
  .I1(mux_o_566),
  .S0(dff_q_6)
);
MUX2 mux_inst_572 (
  .O(mux_o_572),
  .I0(mux_o_568),
  .I1(mux_o_569),
  .S0(dff_q_5)
);
MUX2 mux_inst_573 (
  .O(mux_o_573),
  .I0(mux_o_570),
  .I1(mux_o_567),
  .S0(dff_q_5)
);
MUX2 mux_inst_574 (
  .O(doutb[10]),
  .I0(mux_o_572),
  .I1(mux_o_573),
  .S0(dff_q_4)
);
MUX2 mux_inst_575 (
  .O(mux_o_575),
  .I0(dpx9b_inst_14_doutb[11]),
  .I1(dpx9b_inst_15_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_576 (
  .O(mux_o_576),
  .I0(dpx9b_inst_16_doutb[11]),
  .I1(dpx9b_inst_17_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_577 (
  .O(mux_o_577),
  .I0(dpx9b_inst_18_doutb[11]),
  .I1(dpx9b_inst_19_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_578 (
  .O(mux_o_578),
  .I0(dpx9b_inst_20_doutb[11]),
  .I1(dpx9b_inst_21_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(dpx9b_inst_22_doutb[11]),
  .I1(dpx9b_inst_23_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(dpx9b_inst_24_doutb[11]),
  .I1(dpx9b_inst_25_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_581 (
  .O(mux_o_581),
  .I0(dpx9b_inst_26_doutb[11]),
  .I1(dpx9b_inst_27_doutb[11]),
  .S0(dff_q_7)
);
MUX2 mux_inst_582 (
  .O(mux_o_582),
  .I0(mux_o_575),
  .I1(mux_o_576),
  .S0(dff_q_6)
);
MUX2 mux_inst_583 (
  .O(mux_o_583),
  .I0(mux_o_577),
  .I1(mux_o_578),
  .S0(dff_q_6)
);
MUX2 mux_inst_584 (
  .O(mux_o_584),
  .I0(mux_o_579),
  .I1(mux_o_580),
  .S0(dff_q_6)
);
MUX2 mux_inst_586 (
  .O(mux_o_586),
  .I0(mux_o_582),
  .I1(mux_o_583),
  .S0(dff_q_5)
);
MUX2 mux_inst_587 (
  .O(mux_o_587),
  .I0(mux_o_584),
  .I1(mux_o_581),
  .S0(dff_q_5)
);
MUX2 mux_inst_588 (
  .O(doutb[11]),
  .I0(mux_o_586),
  .I1(mux_o_587),
  .S0(dff_q_4)
);
MUX2 mux_inst_589 (
  .O(mux_o_589),
  .I0(dpx9b_inst_14_doutb[12]),
  .I1(dpx9b_inst_15_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_590 (
  .O(mux_o_590),
  .I0(dpx9b_inst_16_doutb[12]),
  .I1(dpx9b_inst_17_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_591 (
  .O(mux_o_591),
  .I0(dpx9b_inst_18_doutb[12]),
  .I1(dpx9b_inst_19_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_592 (
  .O(mux_o_592),
  .I0(dpx9b_inst_20_doutb[12]),
  .I1(dpx9b_inst_21_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_593 (
  .O(mux_o_593),
  .I0(dpx9b_inst_22_doutb[12]),
  .I1(dpx9b_inst_23_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_594 (
  .O(mux_o_594),
  .I0(dpx9b_inst_24_doutb[12]),
  .I1(dpx9b_inst_25_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_595 (
  .O(mux_o_595),
  .I0(dpx9b_inst_26_doutb[12]),
  .I1(dpx9b_inst_27_doutb[12]),
  .S0(dff_q_7)
);
MUX2 mux_inst_596 (
  .O(mux_o_596),
  .I0(mux_o_589),
  .I1(mux_o_590),
  .S0(dff_q_6)
);
MUX2 mux_inst_597 (
  .O(mux_o_597),
  .I0(mux_o_591),
  .I1(mux_o_592),
  .S0(dff_q_6)
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(mux_o_593),
  .I1(mux_o_594),
  .S0(dff_q_6)
);
MUX2 mux_inst_600 (
  .O(mux_o_600),
  .I0(mux_o_596),
  .I1(mux_o_597),
  .S0(dff_q_5)
);
MUX2 mux_inst_601 (
  .O(mux_o_601),
  .I0(mux_o_598),
  .I1(mux_o_595),
  .S0(dff_q_5)
);
MUX2 mux_inst_602 (
  .O(doutb[12]),
  .I0(mux_o_600),
  .I1(mux_o_601),
  .S0(dff_q_4)
);
MUX2 mux_inst_603 (
  .O(mux_o_603),
  .I0(dpx9b_inst_14_doutb[13]),
  .I1(dpx9b_inst_15_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_604 (
  .O(mux_o_604),
  .I0(dpx9b_inst_16_doutb[13]),
  .I1(dpx9b_inst_17_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_605 (
  .O(mux_o_605),
  .I0(dpx9b_inst_18_doutb[13]),
  .I1(dpx9b_inst_19_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_606 (
  .O(mux_o_606),
  .I0(dpx9b_inst_20_doutb[13]),
  .I1(dpx9b_inst_21_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_607 (
  .O(mux_o_607),
  .I0(dpx9b_inst_22_doutb[13]),
  .I1(dpx9b_inst_23_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_608 (
  .O(mux_o_608),
  .I0(dpx9b_inst_24_doutb[13]),
  .I1(dpx9b_inst_25_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_609 (
  .O(mux_o_609),
  .I0(dpx9b_inst_26_doutb[13]),
  .I1(dpx9b_inst_27_doutb[13]),
  .S0(dff_q_7)
);
MUX2 mux_inst_610 (
  .O(mux_o_610),
  .I0(mux_o_603),
  .I1(mux_o_604),
  .S0(dff_q_6)
);
MUX2 mux_inst_611 (
  .O(mux_o_611),
  .I0(mux_o_605),
  .I1(mux_o_606),
  .S0(dff_q_6)
);
MUX2 mux_inst_612 (
  .O(mux_o_612),
  .I0(mux_o_607),
  .I1(mux_o_608),
  .S0(dff_q_6)
);
MUX2 mux_inst_614 (
  .O(mux_o_614),
  .I0(mux_o_610),
  .I1(mux_o_611),
  .S0(dff_q_5)
);
MUX2 mux_inst_615 (
  .O(mux_o_615),
  .I0(mux_o_612),
  .I1(mux_o_609),
  .S0(dff_q_5)
);
MUX2 mux_inst_616 (
  .O(doutb[13]),
  .I0(mux_o_614),
  .I1(mux_o_615),
  .S0(dff_q_4)
);
MUX2 mux_inst_617 (
  .O(mux_o_617),
  .I0(dpx9b_inst_14_doutb[14]),
  .I1(dpx9b_inst_15_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_618 (
  .O(mux_o_618),
  .I0(dpx9b_inst_16_doutb[14]),
  .I1(dpx9b_inst_17_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_619 (
  .O(mux_o_619),
  .I0(dpx9b_inst_18_doutb[14]),
  .I1(dpx9b_inst_19_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_620 (
  .O(mux_o_620),
  .I0(dpx9b_inst_20_doutb[14]),
  .I1(dpx9b_inst_21_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_621 (
  .O(mux_o_621),
  .I0(dpx9b_inst_22_doutb[14]),
  .I1(dpx9b_inst_23_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_622 (
  .O(mux_o_622),
  .I0(dpx9b_inst_24_doutb[14]),
  .I1(dpx9b_inst_25_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_623 (
  .O(mux_o_623),
  .I0(dpx9b_inst_26_doutb[14]),
  .I1(dpx9b_inst_27_doutb[14]),
  .S0(dff_q_7)
);
MUX2 mux_inst_624 (
  .O(mux_o_624),
  .I0(mux_o_617),
  .I1(mux_o_618),
  .S0(dff_q_6)
);
MUX2 mux_inst_625 (
  .O(mux_o_625),
  .I0(mux_o_619),
  .I1(mux_o_620),
  .S0(dff_q_6)
);
MUX2 mux_inst_626 (
  .O(mux_o_626),
  .I0(mux_o_621),
  .I1(mux_o_622),
  .S0(dff_q_6)
);
MUX2 mux_inst_628 (
  .O(mux_o_628),
  .I0(mux_o_624),
  .I1(mux_o_625),
  .S0(dff_q_5)
);
MUX2 mux_inst_629 (
  .O(mux_o_629),
  .I0(mux_o_626),
  .I1(mux_o_623),
  .S0(dff_q_5)
);
MUX2 mux_inst_630 (
  .O(doutb[14]),
  .I0(mux_o_628),
  .I1(mux_o_629),
  .S0(dff_q_4)
);
MUX2 mux_inst_631 (
  .O(mux_o_631),
  .I0(dpx9b_inst_14_doutb[15]),
  .I1(dpx9b_inst_15_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_632 (
  .O(mux_o_632),
  .I0(dpx9b_inst_16_doutb[15]),
  .I1(dpx9b_inst_17_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_633 (
  .O(mux_o_633),
  .I0(dpx9b_inst_18_doutb[15]),
  .I1(dpx9b_inst_19_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_634 (
  .O(mux_o_634),
  .I0(dpx9b_inst_20_doutb[15]),
  .I1(dpx9b_inst_21_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_635 (
  .O(mux_o_635),
  .I0(dpx9b_inst_22_doutb[15]),
  .I1(dpx9b_inst_23_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_636 (
  .O(mux_o_636),
  .I0(dpx9b_inst_24_doutb[15]),
  .I1(dpx9b_inst_25_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_637 (
  .O(mux_o_637),
  .I0(dpx9b_inst_26_doutb[15]),
  .I1(dpx9b_inst_27_doutb[15]),
  .S0(dff_q_7)
);
MUX2 mux_inst_638 (
  .O(mux_o_638),
  .I0(mux_o_631),
  .I1(mux_o_632),
  .S0(dff_q_6)
);
MUX2 mux_inst_639 (
  .O(mux_o_639),
  .I0(mux_o_633),
  .I1(mux_o_634),
  .S0(dff_q_6)
);
MUX2 mux_inst_640 (
  .O(mux_o_640),
  .I0(mux_o_635),
  .I1(mux_o_636),
  .S0(dff_q_6)
);
MUX2 mux_inst_642 (
  .O(mux_o_642),
  .I0(mux_o_638),
  .I1(mux_o_639),
  .S0(dff_q_5)
);
MUX2 mux_inst_643 (
  .O(mux_o_643),
  .I0(mux_o_640),
  .I1(mux_o_637),
  .S0(dff_q_5)
);
MUX2 mux_inst_644 (
  .O(doutb[15]),
  .I0(mux_o_642),
  .I1(mux_o_643),
  .S0(dff_q_4)
);
MUX2 mux_inst_645 (
  .O(mux_o_645),
  .I0(dpx9b_inst_14_doutb[16]),
  .I1(dpx9b_inst_15_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_646 (
  .O(mux_o_646),
  .I0(dpx9b_inst_16_doutb[16]),
  .I1(dpx9b_inst_17_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_647 (
  .O(mux_o_647),
  .I0(dpx9b_inst_18_doutb[16]),
  .I1(dpx9b_inst_19_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_648 (
  .O(mux_o_648),
  .I0(dpx9b_inst_20_doutb[16]),
  .I1(dpx9b_inst_21_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_649 (
  .O(mux_o_649),
  .I0(dpx9b_inst_22_doutb[16]),
  .I1(dpx9b_inst_23_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_650 (
  .O(mux_o_650),
  .I0(dpx9b_inst_24_doutb[16]),
  .I1(dpx9b_inst_25_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_651 (
  .O(mux_o_651),
  .I0(dpx9b_inst_26_doutb[16]),
  .I1(dpx9b_inst_27_doutb[16]),
  .S0(dff_q_7)
);
MUX2 mux_inst_652 (
  .O(mux_o_652),
  .I0(mux_o_645),
  .I1(mux_o_646),
  .S0(dff_q_6)
);
MUX2 mux_inst_653 (
  .O(mux_o_653),
  .I0(mux_o_647),
  .I1(mux_o_648),
  .S0(dff_q_6)
);
MUX2 mux_inst_654 (
  .O(mux_o_654),
  .I0(mux_o_649),
  .I1(mux_o_650),
  .S0(dff_q_6)
);
MUX2 mux_inst_656 (
  .O(mux_o_656),
  .I0(mux_o_652),
  .I1(mux_o_653),
  .S0(dff_q_5)
);
MUX2 mux_inst_657 (
  .O(mux_o_657),
  .I0(mux_o_654),
  .I1(mux_o_651),
  .S0(dff_q_5)
);
MUX2 mux_inst_658 (
  .O(doutb[16]),
  .I0(mux_o_656),
  .I1(mux_o_657),
  .S0(dff_q_4)
);
MUX2 mux_inst_659 (
  .O(mux_o_659),
  .I0(dpx9b_inst_14_doutb[17]),
  .I1(dpx9b_inst_15_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_660 (
  .O(mux_o_660),
  .I0(dpx9b_inst_16_doutb[17]),
  .I1(dpx9b_inst_17_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_661 (
  .O(mux_o_661),
  .I0(dpx9b_inst_18_doutb[17]),
  .I1(dpx9b_inst_19_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_662 (
  .O(mux_o_662),
  .I0(dpx9b_inst_20_doutb[17]),
  .I1(dpx9b_inst_21_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_663 (
  .O(mux_o_663),
  .I0(dpx9b_inst_22_doutb[17]),
  .I1(dpx9b_inst_23_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_664 (
  .O(mux_o_664),
  .I0(dpx9b_inst_24_doutb[17]),
  .I1(dpx9b_inst_25_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_665 (
  .O(mux_o_665),
  .I0(dpx9b_inst_26_doutb[17]),
  .I1(dpx9b_inst_27_doutb[17]),
  .S0(dff_q_7)
);
MUX2 mux_inst_666 (
  .O(mux_o_666),
  .I0(mux_o_659),
  .I1(mux_o_660),
  .S0(dff_q_6)
);
MUX2 mux_inst_667 (
  .O(mux_o_667),
  .I0(mux_o_661),
  .I1(mux_o_662),
  .S0(dff_q_6)
);
MUX2 mux_inst_668 (
  .O(mux_o_668),
  .I0(mux_o_663),
  .I1(mux_o_664),
  .S0(dff_q_6)
);
MUX2 mux_inst_670 (
  .O(mux_o_670),
  .I0(mux_o_666),
  .I1(mux_o_667),
  .S0(dff_q_5)
);
MUX2 mux_inst_671 (
  .O(mux_o_671),
  .I0(mux_o_668),
  .I1(mux_o_665),
  .S0(dff_q_5)
);
MUX2 mux_inst_672 (
  .O(doutb[17]),
  .I0(mux_o_670),
  .I1(mux_o_671),
  .S0(dff_q_4)
);
MUX2 mux_inst_673 (
  .O(mux_o_673),
  .I0(dpx9b_inst_28_doutb[18]),
  .I1(dpx9b_inst_29_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_674 (
  .O(mux_o_674),
  .I0(dpx9b_inst_30_doutb[18]),
  .I1(dpx9b_inst_31_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_675 (
  .O(mux_o_675),
  .I0(dpx9b_inst_32_doutb[18]),
  .I1(dpx9b_inst_33_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_676 (
  .O(mux_o_676),
  .I0(dpx9b_inst_34_doutb[18]),
  .I1(dpx9b_inst_35_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_677 (
  .O(mux_o_677),
  .I0(dpx9b_inst_36_doutb[18]),
  .I1(dpx9b_inst_37_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_678 (
  .O(mux_o_678),
  .I0(dpx9b_inst_38_doutb[18]),
  .I1(dpx9b_inst_39_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_679 (
  .O(mux_o_679),
  .I0(dpx9b_inst_40_doutb[18]),
  .I1(dpx9b_inst_41_doutb[18]),
  .S0(dff_q_7)
);
MUX2 mux_inst_680 (
  .O(mux_o_680),
  .I0(mux_o_673),
  .I1(mux_o_674),
  .S0(dff_q_6)
);
MUX2 mux_inst_681 (
  .O(mux_o_681),
  .I0(mux_o_675),
  .I1(mux_o_676),
  .S0(dff_q_6)
);
MUX2 mux_inst_682 (
  .O(mux_o_682),
  .I0(mux_o_677),
  .I1(mux_o_678),
  .S0(dff_q_6)
);
MUX2 mux_inst_684 (
  .O(mux_o_684),
  .I0(mux_o_680),
  .I1(mux_o_681),
  .S0(dff_q_5)
);
MUX2 mux_inst_685 (
  .O(mux_o_685),
  .I0(mux_o_682),
  .I1(mux_o_679),
  .S0(dff_q_5)
);
MUX2 mux_inst_686 (
  .O(doutb[18]),
  .I0(mux_o_684),
  .I1(mux_o_685),
  .S0(dff_q_4)
);
MUX2 mux_inst_687 (
  .O(mux_o_687),
  .I0(dpx9b_inst_28_doutb[19]),
  .I1(dpx9b_inst_29_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_688 (
  .O(mux_o_688),
  .I0(dpx9b_inst_30_doutb[19]),
  .I1(dpx9b_inst_31_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_689 (
  .O(mux_o_689),
  .I0(dpx9b_inst_32_doutb[19]),
  .I1(dpx9b_inst_33_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_690 (
  .O(mux_o_690),
  .I0(dpx9b_inst_34_doutb[19]),
  .I1(dpx9b_inst_35_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_691 (
  .O(mux_o_691),
  .I0(dpx9b_inst_36_doutb[19]),
  .I1(dpx9b_inst_37_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_692 (
  .O(mux_o_692),
  .I0(dpx9b_inst_38_doutb[19]),
  .I1(dpx9b_inst_39_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_693 (
  .O(mux_o_693),
  .I0(dpx9b_inst_40_doutb[19]),
  .I1(dpx9b_inst_41_doutb[19]),
  .S0(dff_q_7)
);
MUX2 mux_inst_694 (
  .O(mux_o_694),
  .I0(mux_o_687),
  .I1(mux_o_688),
  .S0(dff_q_6)
);
MUX2 mux_inst_695 (
  .O(mux_o_695),
  .I0(mux_o_689),
  .I1(mux_o_690),
  .S0(dff_q_6)
);
MUX2 mux_inst_696 (
  .O(mux_o_696),
  .I0(mux_o_691),
  .I1(mux_o_692),
  .S0(dff_q_6)
);
MUX2 mux_inst_698 (
  .O(mux_o_698),
  .I0(mux_o_694),
  .I1(mux_o_695),
  .S0(dff_q_5)
);
MUX2 mux_inst_699 (
  .O(mux_o_699),
  .I0(mux_o_696),
  .I1(mux_o_693),
  .S0(dff_q_5)
);
MUX2 mux_inst_700 (
  .O(doutb[19]),
  .I0(mux_o_698),
  .I1(mux_o_699),
  .S0(dff_q_4)
);
MUX2 mux_inst_701 (
  .O(mux_o_701),
  .I0(dpx9b_inst_28_doutb[20]),
  .I1(dpx9b_inst_29_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_702 (
  .O(mux_o_702),
  .I0(dpx9b_inst_30_doutb[20]),
  .I1(dpx9b_inst_31_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_703 (
  .O(mux_o_703),
  .I0(dpx9b_inst_32_doutb[20]),
  .I1(dpx9b_inst_33_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_704 (
  .O(mux_o_704),
  .I0(dpx9b_inst_34_doutb[20]),
  .I1(dpx9b_inst_35_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_705 (
  .O(mux_o_705),
  .I0(dpx9b_inst_36_doutb[20]),
  .I1(dpx9b_inst_37_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_706 (
  .O(mux_o_706),
  .I0(dpx9b_inst_38_doutb[20]),
  .I1(dpx9b_inst_39_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_707 (
  .O(mux_o_707),
  .I0(dpx9b_inst_40_doutb[20]),
  .I1(dpx9b_inst_41_doutb[20]),
  .S0(dff_q_7)
);
MUX2 mux_inst_708 (
  .O(mux_o_708),
  .I0(mux_o_701),
  .I1(mux_o_702),
  .S0(dff_q_6)
);
MUX2 mux_inst_709 (
  .O(mux_o_709),
  .I0(mux_o_703),
  .I1(mux_o_704),
  .S0(dff_q_6)
);
MUX2 mux_inst_710 (
  .O(mux_o_710),
  .I0(mux_o_705),
  .I1(mux_o_706),
  .S0(dff_q_6)
);
MUX2 mux_inst_712 (
  .O(mux_o_712),
  .I0(mux_o_708),
  .I1(mux_o_709),
  .S0(dff_q_5)
);
MUX2 mux_inst_713 (
  .O(mux_o_713),
  .I0(mux_o_710),
  .I1(mux_o_707),
  .S0(dff_q_5)
);
MUX2 mux_inst_714 (
  .O(doutb[20]),
  .I0(mux_o_712),
  .I1(mux_o_713),
  .S0(dff_q_4)
);
MUX2 mux_inst_715 (
  .O(mux_o_715),
  .I0(dpx9b_inst_28_doutb[21]),
  .I1(dpx9b_inst_29_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_716 (
  .O(mux_o_716),
  .I0(dpx9b_inst_30_doutb[21]),
  .I1(dpx9b_inst_31_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_717 (
  .O(mux_o_717),
  .I0(dpx9b_inst_32_doutb[21]),
  .I1(dpx9b_inst_33_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_718 (
  .O(mux_o_718),
  .I0(dpx9b_inst_34_doutb[21]),
  .I1(dpx9b_inst_35_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_719 (
  .O(mux_o_719),
  .I0(dpx9b_inst_36_doutb[21]),
  .I1(dpx9b_inst_37_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_720 (
  .O(mux_o_720),
  .I0(dpx9b_inst_38_doutb[21]),
  .I1(dpx9b_inst_39_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_721 (
  .O(mux_o_721),
  .I0(dpx9b_inst_40_doutb[21]),
  .I1(dpx9b_inst_41_doutb[21]),
  .S0(dff_q_7)
);
MUX2 mux_inst_722 (
  .O(mux_o_722),
  .I0(mux_o_715),
  .I1(mux_o_716),
  .S0(dff_q_6)
);
MUX2 mux_inst_723 (
  .O(mux_o_723),
  .I0(mux_o_717),
  .I1(mux_o_718),
  .S0(dff_q_6)
);
MUX2 mux_inst_724 (
  .O(mux_o_724),
  .I0(mux_o_719),
  .I1(mux_o_720),
  .S0(dff_q_6)
);
MUX2 mux_inst_726 (
  .O(mux_o_726),
  .I0(mux_o_722),
  .I1(mux_o_723),
  .S0(dff_q_5)
);
MUX2 mux_inst_727 (
  .O(mux_o_727),
  .I0(mux_o_724),
  .I1(mux_o_721),
  .S0(dff_q_5)
);
MUX2 mux_inst_728 (
  .O(doutb[21]),
  .I0(mux_o_726),
  .I1(mux_o_727),
  .S0(dff_q_4)
);
MUX2 mux_inst_729 (
  .O(mux_o_729),
  .I0(dpx9b_inst_28_doutb[22]),
  .I1(dpx9b_inst_29_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_730 (
  .O(mux_o_730),
  .I0(dpx9b_inst_30_doutb[22]),
  .I1(dpx9b_inst_31_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_731 (
  .O(mux_o_731),
  .I0(dpx9b_inst_32_doutb[22]),
  .I1(dpx9b_inst_33_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_732 (
  .O(mux_o_732),
  .I0(dpx9b_inst_34_doutb[22]),
  .I1(dpx9b_inst_35_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_733 (
  .O(mux_o_733),
  .I0(dpx9b_inst_36_doutb[22]),
  .I1(dpx9b_inst_37_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_734 (
  .O(mux_o_734),
  .I0(dpx9b_inst_38_doutb[22]),
  .I1(dpx9b_inst_39_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_735 (
  .O(mux_o_735),
  .I0(dpx9b_inst_40_doutb[22]),
  .I1(dpx9b_inst_41_doutb[22]),
  .S0(dff_q_7)
);
MUX2 mux_inst_736 (
  .O(mux_o_736),
  .I0(mux_o_729),
  .I1(mux_o_730),
  .S0(dff_q_6)
);
MUX2 mux_inst_737 (
  .O(mux_o_737),
  .I0(mux_o_731),
  .I1(mux_o_732),
  .S0(dff_q_6)
);
MUX2 mux_inst_738 (
  .O(mux_o_738),
  .I0(mux_o_733),
  .I1(mux_o_734),
  .S0(dff_q_6)
);
MUX2 mux_inst_740 (
  .O(mux_o_740),
  .I0(mux_o_736),
  .I1(mux_o_737),
  .S0(dff_q_5)
);
MUX2 mux_inst_741 (
  .O(mux_o_741),
  .I0(mux_o_738),
  .I1(mux_o_735),
  .S0(dff_q_5)
);
MUX2 mux_inst_742 (
  .O(doutb[22]),
  .I0(mux_o_740),
  .I1(mux_o_741),
  .S0(dff_q_4)
);
MUX2 mux_inst_743 (
  .O(mux_o_743),
  .I0(dpx9b_inst_28_doutb[23]),
  .I1(dpx9b_inst_29_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_744 (
  .O(mux_o_744),
  .I0(dpx9b_inst_30_doutb[23]),
  .I1(dpx9b_inst_31_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_745 (
  .O(mux_o_745),
  .I0(dpx9b_inst_32_doutb[23]),
  .I1(dpx9b_inst_33_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_746 (
  .O(mux_o_746),
  .I0(dpx9b_inst_34_doutb[23]),
  .I1(dpx9b_inst_35_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_747 (
  .O(mux_o_747),
  .I0(dpx9b_inst_36_doutb[23]),
  .I1(dpx9b_inst_37_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_748 (
  .O(mux_o_748),
  .I0(dpx9b_inst_38_doutb[23]),
  .I1(dpx9b_inst_39_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_749 (
  .O(mux_o_749),
  .I0(dpx9b_inst_40_doutb[23]),
  .I1(dpx9b_inst_41_doutb[23]),
  .S0(dff_q_7)
);
MUX2 mux_inst_750 (
  .O(mux_o_750),
  .I0(mux_o_743),
  .I1(mux_o_744),
  .S0(dff_q_6)
);
MUX2 mux_inst_751 (
  .O(mux_o_751),
  .I0(mux_o_745),
  .I1(mux_o_746),
  .S0(dff_q_6)
);
MUX2 mux_inst_752 (
  .O(mux_o_752),
  .I0(mux_o_747),
  .I1(mux_o_748),
  .S0(dff_q_6)
);
MUX2 mux_inst_754 (
  .O(mux_o_754),
  .I0(mux_o_750),
  .I1(mux_o_751),
  .S0(dff_q_5)
);
MUX2 mux_inst_755 (
  .O(mux_o_755),
  .I0(mux_o_752),
  .I1(mux_o_749),
  .S0(dff_q_5)
);
MUX2 mux_inst_756 (
  .O(doutb[23]),
  .I0(mux_o_754),
  .I1(mux_o_755),
  .S0(dff_q_4)
);
MUX2 mux_inst_757 (
  .O(mux_o_757),
  .I0(dpx9b_inst_28_doutb[24]),
  .I1(dpx9b_inst_29_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_758 (
  .O(mux_o_758),
  .I0(dpx9b_inst_30_doutb[24]),
  .I1(dpx9b_inst_31_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_759 (
  .O(mux_o_759),
  .I0(dpx9b_inst_32_doutb[24]),
  .I1(dpx9b_inst_33_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_760 (
  .O(mux_o_760),
  .I0(dpx9b_inst_34_doutb[24]),
  .I1(dpx9b_inst_35_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_761 (
  .O(mux_o_761),
  .I0(dpx9b_inst_36_doutb[24]),
  .I1(dpx9b_inst_37_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_762 (
  .O(mux_o_762),
  .I0(dpx9b_inst_38_doutb[24]),
  .I1(dpx9b_inst_39_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_763 (
  .O(mux_o_763),
  .I0(dpx9b_inst_40_doutb[24]),
  .I1(dpx9b_inst_41_doutb[24]),
  .S0(dff_q_7)
);
MUX2 mux_inst_764 (
  .O(mux_o_764),
  .I0(mux_o_757),
  .I1(mux_o_758),
  .S0(dff_q_6)
);
MUX2 mux_inst_765 (
  .O(mux_o_765),
  .I0(mux_o_759),
  .I1(mux_o_760),
  .S0(dff_q_6)
);
MUX2 mux_inst_766 (
  .O(mux_o_766),
  .I0(mux_o_761),
  .I1(mux_o_762),
  .S0(dff_q_6)
);
MUX2 mux_inst_768 (
  .O(mux_o_768),
  .I0(mux_o_764),
  .I1(mux_o_765),
  .S0(dff_q_5)
);
MUX2 mux_inst_769 (
  .O(mux_o_769),
  .I0(mux_o_766),
  .I1(mux_o_763),
  .S0(dff_q_5)
);
MUX2 mux_inst_770 (
  .O(doutb[24]),
  .I0(mux_o_768),
  .I1(mux_o_769),
  .S0(dff_q_4)
);
MUX2 mux_inst_771 (
  .O(mux_o_771),
  .I0(dpx9b_inst_28_doutb[25]),
  .I1(dpx9b_inst_29_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_772 (
  .O(mux_o_772),
  .I0(dpx9b_inst_30_doutb[25]),
  .I1(dpx9b_inst_31_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_773 (
  .O(mux_o_773),
  .I0(dpx9b_inst_32_doutb[25]),
  .I1(dpx9b_inst_33_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_774 (
  .O(mux_o_774),
  .I0(dpx9b_inst_34_doutb[25]),
  .I1(dpx9b_inst_35_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_775 (
  .O(mux_o_775),
  .I0(dpx9b_inst_36_doutb[25]),
  .I1(dpx9b_inst_37_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_776 (
  .O(mux_o_776),
  .I0(dpx9b_inst_38_doutb[25]),
  .I1(dpx9b_inst_39_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_777 (
  .O(mux_o_777),
  .I0(dpx9b_inst_40_doutb[25]),
  .I1(dpx9b_inst_41_doutb[25]),
  .S0(dff_q_7)
);
MUX2 mux_inst_778 (
  .O(mux_o_778),
  .I0(mux_o_771),
  .I1(mux_o_772),
  .S0(dff_q_6)
);
MUX2 mux_inst_779 (
  .O(mux_o_779),
  .I0(mux_o_773),
  .I1(mux_o_774),
  .S0(dff_q_6)
);
MUX2 mux_inst_780 (
  .O(mux_o_780),
  .I0(mux_o_775),
  .I1(mux_o_776),
  .S0(dff_q_6)
);
MUX2 mux_inst_782 (
  .O(mux_o_782),
  .I0(mux_o_778),
  .I1(mux_o_779),
  .S0(dff_q_5)
);
MUX2 mux_inst_783 (
  .O(mux_o_783),
  .I0(mux_o_780),
  .I1(mux_o_777),
  .S0(dff_q_5)
);
MUX2 mux_inst_784 (
  .O(doutb[25]),
  .I0(mux_o_782),
  .I1(mux_o_783),
  .S0(dff_q_4)
);
MUX2 mux_inst_785 (
  .O(mux_o_785),
  .I0(dpx9b_inst_28_doutb[26]),
  .I1(dpx9b_inst_29_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_786 (
  .O(mux_o_786),
  .I0(dpx9b_inst_30_doutb[26]),
  .I1(dpx9b_inst_31_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_787 (
  .O(mux_o_787),
  .I0(dpx9b_inst_32_doutb[26]),
  .I1(dpx9b_inst_33_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_788 (
  .O(mux_o_788),
  .I0(dpx9b_inst_34_doutb[26]),
  .I1(dpx9b_inst_35_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_789 (
  .O(mux_o_789),
  .I0(dpx9b_inst_36_doutb[26]),
  .I1(dpx9b_inst_37_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_790 (
  .O(mux_o_790),
  .I0(dpx9b_inst_38_doutb[26]),
  .I1(dpx9b_inst_39_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_791 (
  .O(mux_o_791),
  .I0(dpx9b_inst_40_doutb[26]),
  .I1(dpx9b_inst_41_doutb[26]),
  .S0(dff_q_7)
);
MUX2 mux_inst_792 (
  .O(mux_o_792),
  .I0(mux_o_785),
  .I1(mux_o_786),
  .S0(dff_q_6)
);
MUX2 mux_inst_793 (
  .O(mux_o_793),
  .I0(mux_o_787),
  .I1(mux_o_788),
  .S0(dff_q_6)
);
MUX2 mux_inst_794 (
  .O(mux_o_794),
  .I0(mux_o_789),
  .I1(mux_o_790),
  .S0(dff_q_6)
);
MUX2 mux_inst_796 (
  .O(mux_o_796),
  .I0(mux_o_792),
  .I1(mux_o_793),
  .S0(dff_q_5)
);
MUX2 mux_inst_797 (
  .O(mux_o_797),
  .I0(mux_o_794),
  .I1(mux_o_791),
  .S0(dff_q_5)
);
MUX2 mux_inst_798 (
  .O(doutb[26]),
  .I0(mux_o_796),
  .I1(mux_o_797),
  .S0(dff_q_4)
);
MUX2 mux_inst_806 (
  .O(mux_o_806),
  .I0(dpb_inst_46_doutb[27]),
  .I1(dpb_inst_48_doutb[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_807 (
  .O(doutb[27]),
  .I0(dpb_inst_42_doutb[27]),
  .I1(mux_o_806),
  .S0(dff_q_4)
);
MUX2 mux_inst_815 (
  .O(mux_o_815),
  .I0(dpb_inst_46_doutb[28]),
  .I1(dpb_inst_48_doutb[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_816 (
  .O(doutb[28]),
  .I0(dpb_inst_43_doutb[28]),
  .I1(mux_o_815),
  .S0(dff_q_4)
);
MUX2 mux_inst_824 (
  .O(mux_o_824),
  .I0(dpb_inst_47_doutb[29]),
  .I1(dpb_inst_48_doutb[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_825 (
  .O(doutb[29]),
  .I0(dpb_inst_44_doutb[29]),
  .I1(mux_o_824),
  .S0(dff_q_4)
);
MUX2 mux_inst_833 (
  .O(mux_o_833),
  .I0(dpb_inst_47_doutb[30]),
  .I1(dpb_inst_48_doutb[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_834 (
  .O(doutb[30]),
  .I0(dpb_inst_45_doutb[30]),
  .I1(mux_o_833),
  .S0(dff_q_4)
);
MUX2 mux_inst_841 (
  .O(doutb[31]),
  .I0(dpb_inst_49_doutb[31]),
  .I1(dpb_inst_50_doutb[31]),
  .S0(dff_q_4)
);
endmodule //Gowin_DPB
